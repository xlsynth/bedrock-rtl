// Copyright 2024 The Bedrock-RTL Authors
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//     http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.

// Bridge AXI4-Lite to APB Bridge
//
// Converts an AXI4-Lite interface to an APB interface.

`include "br_asserts_internal.svh"
`include "br_registers.svh"

module br_amba_axil2apb #(
    parameter int AddrWidth = 40,
    parameter int DataWidth = 64
) (
    input clk,
    input rst,  // Synchronous, active-high reset

    // AXI4-Lite interface
    input  logic [    AddrWidth-1:0] awaddr,
    input  logic [              2:0] awprot,
    input  logic                     awvalid,
    output logic                     awready,
    input  logic [    DataWidth-1:0] wdata,
    input  logic [(DataWidth/8)-1:0] wstrb,
    input  logic                     wvalid,
    output logic                     wready,
    output logic [              1:0] bresp,
    output logic                     bvalid,
    input  logic                     bready,
    input  logic [    AddrWidth-1:0] araddr,
    input  logic [              2:0] arprot,
    input  logic                     arvalid,
    output logic                     arready,
    output logic [    DataWidth-1:0] rdata,
    output logic [              1:0] rresp,
    output logic                     rvalid,
    input  logic                     rready,

    // APB interface
    output logic [    AddrWidth-1:0] paddr,
    output logic                     psel,
    output logic                     penable,
    output logic [              2:0] pprot,
    output logic [(DataWidth/8)-1:0] pstrb,
    output logic                     pwrite,
    output logic [    DataWidth-1:0] pwdata,
    input  logic [    DataWidth-1:0] prdata,
    input  logic                     pready,
    input  logic                     pslverr
);

  typedef enum logic [3:0] {
    IDLE   = 4'b0001,
    SETUP  = 4'b0010,
    ACCESS = 4'b0100,
    RESP   = 4'b1000
  } apb_state_t;
  apb_state_t apb_state, apb_state_next;

  logic [AddrWidth-1:0] addr_reg, addr_next;
  logic [DataWidth-1:0] data_reg;
  logic [(DataWidth/8)-1:0] strb_reg;
  logic [2:0] prot_reg, prot_next;
  logic resp_reg;
  logic write_reg;
  logic arb_write_req, arb_write_grant;
  logic arb_read_req, arb_read_grant;
  logic arb_any_grant;
  logic write_txn, write_txn_next;
  logic read_txn, read_txn_next;
  logic write_done, write_done_next;
  logic read_done, read_done_next;

  `BR_REGLN(addr_reg, addr_next, arb_any_grant)
  `BR_REGLN(data_reg, wdata, arb_any_grant)
  `BR_REGLN(write_reg, write_txn, arb_any_grant)
  `BR_REGLN(strb_reg, wstrb, arb_any_grant)
  `BR_REGLN(prot_reg, prot_next, arb_any_grant)
  `BR_REGLN(resp_reg, pslverr, (apb_state == ACCESS) && pready)
  `BR_REGLN(rdata, prdata, read_done)
  `BR_REG(write_txn, write_txn_next)
  `BR_REG(read_txn, read_txn_next)
  `BR_REG(write_done, write_done_next)
  `BR_REG(read_done, read_done_next)
  `BR_REGI(apb_state, apb_state_next, IDLE)

  // Arbitrate between read and write transactions
  br_arb_rr #(
      .NumRequesters(2)
  ) br_arb_rr (
      .clk(clk),
      .rst(rst),
      .enable_priority_update(1'b0),
      .request({arb_write_req, arb_read_req}),
      .grant({arb_write_grant, arb_read_grant})
  );

  // Arbiter request signals
  assign arb_write_req = awvalid && wvalid && ~bvalid && (apb_state == IDLE);
  assign arb_read_req = arvalid && ~rvalid && (apb_state == IDLE);
  assign arb_any_grant = arb_write_grant || arb_read_grant;

  // Save the address and data for the transaction
  assign addr_next = arb_write_grant ? awaddr : araddr;
  assign prot_next = arb_write_grant ? awprot : arprot;

  // Track transaction state
  assign write_txn_next = (write_txn && ~write_done) || (~write_txn && arb_write_grant);
  assign read_txn_next = (read_txn && ~read_done) || (~read_txn && arb_read_grant);

  // Track transaction completion
  assign write_done_next = bvalid && bready;
  assign read_done_next = rvalid && rready;

  // APB state machine
  // ri lint_check_off GRAY_CODE_FSM
  always_comb begin
    // Default next state
    apb_state_next = apb_state;

    unique case (apb_state)  // ri lint_check_waive FSM_DEFAULT_REQ
      IDLE: begin
        if (arb_any_grant) begin
          apb_state_next = SETUP;
        end
      end
      SETUP: begin
        apb_state_next = ACCESS;
      end
      ACCESS: begin
        if (pready) begin
          apb_state_next = RESP;
        end
      end
      RESP: begin
        if (write_done_next || read_done_next) begin
          apb_state_next = IDLE;
        end
      end
    endcase
  end
  // ri lint_check_on GRAY_CODE_FSM

  // AXI4-Lite signal generation
  assign awready = arb_write_grant;
  assign wready = arb_write_grant;
  assign bvalid = (apb_state == RESP) && write_txn;
  assign bresp = {resp_reg, 1'b0};  // ri lint_check_waive CONST_ASSIGN CONST_OUTPUT
  assign arready = arb_read_grant;
  assign rvalid = (apb_state == RESP) && read_txn;
  assign rresp = {resp_reg, 1'b0};  // ri lint_check_waive CONST_ASSIGN CONST_OUTPUT

  // APB signal generation
  assign psel = (apb_state != IDLE);
  assign penable = (apb_state == ACCESS);
  assign paddr = addr_reg;
  assign pwdata = data_reg;
  assign pwrite = write_reg;
  assign pprot = prot_reg;
  assign pstrb = strb_reg;

  //------------------------------------------
  // Implementation checks
  //------------------------------------------

  `BR_ASSERT_IMPL(apb_state_next_known_a, !$isunknown(apb_state_next))

endmodule : br_amba_axil2apb
