// Copyright 2024-2025 The Bedrock-RTL Authors
//
// Licensed under the Apache License, Version 2.0 (the "License");
// Copyright 2024-2025 The Bedrock-RTL Authors
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//     http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.


// verilog_format: off
// verilog_lint: waive-start line-length

// Bedrock-RTL Single-Error-Correcting, Double-Error-Detecting (SECDED - Hsiao) Encoder
//
// Encodes a message using a single-error-correcting, double-error-detecting
// linear block code in systematic form (in layperson's terms: a Hsiao SECDED [1] encoder,
// closely related to Hamming codes).
//
// Systematic form means that the codeword is formed by appending the
// calculated parity bits to the message, i.e., the code has the property
// that the message bits are 1:1 with a slice of bits in the codeword (if they
// have not been corrupted).
//
// In Bedrock ECC libs, our convention is to always append the parity bits on
// the MSbs:
//     codeword == {parity, message}
//
// This module has parameterizable latency. By default, it is purely combinational,
// but it can have up to 2 cycles of delay (RegisterInputs and RegisterOutputs).
// The initiation interval is always 1 cycle.
//
// Any data width >= 4 is supported, up to a maximum of 1024. It is internally zero-padded up to
// the largest message width supported by the number of parity bits before being encoded.
// The following table outlines the number of parity bits required for different message widths.
//
// | Message Width (k) | Parity Width (r) | Codeword Width (n)|
// |-------------------|------------------|-------------------|
// | 4                 | 4                | 8                 |
// | 11                | 5                | 16                |
// | 26                | 6                | 32                |
// | 57                | 7                | 64                |
// | 120               | 8                | 128               |
// | 247               | 9                | 256               |
// | 502               | 10               | 512               |
// | 1013              | 11               | 1024              |
// | 2036              | 12               | 2048              |
//
// The number of parity bits must be one of the values in the table above
// or the module will not elaborate.
//
// References:
// [1] https://ieeexplore.ieee.org/abstract/document/5391627

`include "br_asserts.svh"
`include "br_asserts_internal.svh"
`include "br_assign.svh"
`include "br_unused.svh"

module br_ecc_secded_encoder #(
    parameter int DataWidth = 4,  // Must be at least 4
    parameter int ParityWidth = 4,  // Must be at least 4 and at most 12
    // If 1, then insert a pipeline register at the input.
    parameter bit RegisterInputs = 0,
    // If 1, then insert a pipeline register at the output.
    parameter bit RegisterOutputs = 0,
    // If 1, then assert there are no valid bits asserted at the end of the test.
    parameter bit EnableAssertFinalNotValid = 1,
    localparam int OutputWidth = DataWidth + ParityWidth,
    localparam int MessageWidth = br_ecc::get_max_message_width(ParityWidth),
    localparam int CodewordWidth = MessageWidth + ParityWidth
) (
    // Positive edge-triggered clock.
    input  logic                     clk,
    // Synchronous active-high reset.
    input  logic                     rst,
    input  logic                     data_valid,
    input  logic [    DataWidth-1:0] data,
    output logic                     enc_valid,
    output logic [    DataWidth-1:0] enc_data,
    output logic [  ParityWidth-1:0] enc_parity,
    // A concatenation of {enc_parity, 0 padding, enc_data}, i.e.,
    // {enc_parity, message}
    output logic [CodewordWidth-1:0] enc_codeword
);

  // ri lint_check_waive PARAM_NOT_USED
  localparam int Latency = RegisterInputs + RegisterOutputs;

  //------------------------------------------
  // Integration checks
  //------------------------------------------
  `BR_ASSERT_STATIC(data_width_gte_4_a, DataWidth >= 4)
  `BR_ASSERT_STATIC(parity_width_gte_4_a, ParityWidth >= 4)
  `BR_ASSERT_STATIC(parity_width_lte_12_a, ParityWidth <= 12)
  `BR_ASSERT_STATIC(codeword_width_pow_of_2_a, br_math::is_power_of_2(CodewordWidth))
  `BR_ASSERT_STATIC(data_width_fits_in_message_width_a, DataWidth <= MessageWidth)
  `BR_ASSERT_STATIC(right_sized_parity_bits_a, DataWidth > br_ecc::get_max_message_width(ParityWidth - 1))

  //------------------------------------------
  // Implementation
  //------------------------------------------

  //------
  // Optionally register the input signals.
  //------
  logic data_valid_d;
  logic [DataWidth-1:0] data_d;

  br_delay_valid #(
      .Width(DataWidth),
      .NumStages(RegisterInputs == 1 ? 1 : 0),
      .EnableAssertFinalNotValid(EnableAssertFinalNotValid)
  ) br_delay_valid_inputs (
      .clk,
      .rst,
      .in_valid(data_valid),
      .in(data),
      .out_valid(data_valid_d),
      .out(data_d),
      .out_valid_stages(),  // unused
      .out_stages()  // unused
  );

  //------
  // Pad the data to the message width.
  //------

  localparam int PadWidth = MessageWidth - DataWidth;
  logic [MessageWidth-1:0] m;

  if (PadWidth > 0) begin : gen_pad
    assign m = { {PadWidth{1'b0} }, data_d};
  end else begin : gen_no_pad
    assign m = data_d;
  end

  //------
  // Compute parity bits.
  //------
  logic [ParityWidth-1:0] parity;

  // ri lint_check_off EXPR_ID_LIMIT

  if ((CodewordWidth == 8) && (MessageWidth == 4)) begin : gen_8_4
    `BR_ASSERT_STATIC(parity_width_matches_a, ParityWidth == 4)
    assign parity[0] = m[1] ^ m[2] ^ m[3];
    assign parity[1] = m[0] ^ m[2] ^ m[3];
    assign parity[2] = m[0] ^ m[1] ^ m[3];
    assign parity[3] = m[0] ^ m[1] ^ m[2];
  end else if ((CodewordWidth == 16) && (MessageWidth == 11)) begin : gen_16_11
    `BR_ASSERT_STATIC(parity_width_matches_a, ParityWidth == 5)
    assign parity[0] = m[0] ^ m[2] ^ m[4] ^ m[5] ^ m[7] ^ m[8] ^ m[10];
    assign parity[1] = m[0] ^ m[2] ^ m[3] ^ m[5] ^ m[6] ^ m[9] ^ m[10];
    assign parity[2] = m[0] ^ m[1] ^ m[3] ^ m[5] ^ m[7] ^ m[8] ^ m[9];
    assign parity[3] = m[0] ^ m[1] ^ m[3] ^ m[4] ^ m[6] ^ m[8] ^ m[10];
    assign parity[4] = m[0] ^ m[1] ^ m[2] ^ m[4] ^ m[6] ^ m[7] ^ m[9];
  end else if ((CodewordWidth == 32) && (MessageWidth == 26)) begin : gen_32_26
    `BR_ASSERT_STATIC(parity_width_matches_a, ParityWidth == 6)
    assign parity[0] = m[1] ^ m[3] ^ m[5] ^ m[6] ^ m[9] ^ m[11] ^ m[12] ^ m[15] ^ m[16] ^ m[18] ^ m[21] ^ m[22] ^ m[23] ^ m[24] ^ m[25];
    assign parity[1] = m[1] ^ m[3] ^ m[4] ^ m[7] ^ m[9] ^ m[10] ^ m[13] ^ m[14] ^ m[17] ^ m[18] ^ m[20] ^ m[22] ^ m[23] ^ m[24] ^ m[25];
    assign parity[2] = m[1] ^ m[2] ^ m[5] ^ m[7] ^ m[8] ^ m[11] ^ m[13] ^ m[14] ^ m[16] ^ m[19] ^ m[20] ^ m[21] ^ m[23] ^ m[24] ^ m[25];
    assign parity[3] = m[0] ^ m[3] ^ m[5] ^ m[7] ^ m[8] ^ m[10] ^ m[12] ^ m[15] ^ m[17] ^ m[19] ^ m[20] ^ m[21] ^ m[22] ^ m[24] ^ m[25];
    assign parity[4] = m[0] ^ m[2] ^ m[4] ^ m[6] ^ m[9] ^ m[11] ^ m[13] ^ m[15] ^ m[17] ^ m[19] ^ m[20] ^ m[21] ^ m[22] ^ m[23] ^ m[25];
    assign parity[5] = m[0] ^ m[2] ^ m[4] ^ m[6] ^ m[8] ^ m[10] ^ m[12] ^ m[14] ^ m[16] ^ m[18] ^ m[20] ^ m[21] ^ m[22] ^ m[23] ^ m[24];
  end else if ((CodewordWidth == 64) && (MessageWidth == 57)) begin : gen_64_57
    `BR_ASSERT_STATIC(parity_width_matches_a, ParityWidth == 7)
    assign parity[0] = m[0] ^ m[2] ^ m[4] ^ m[6] ^ m[8] ^ m[10] ^ m[12] ^ m[14] ^ m[15] ^ m[17] ^ m[20] ^ m[22] ^ m[24] ^ m[26] ^ m[27] ^ m[30] ^ m[32] ^ m[33] ^ m[35] ^ m[38] ^ m[39] ^ m[42] ^ m[44] ^ m[45] ^ m[47] ^ m[48] ^ m[49] ^ m[50] ^ m[52] ^ m[54] ^ m[56];
    assign parity[1] = m[0] ^ m[2] ^ m[4] ^ m[6] ^ m[8] ^ m[10] ^ m[11] ^ m[13] ^ m[16] ^ m[18] ^ m[20] ^ m[22] ^ m[23] ^ m[26] ^ m[28] ^ m[29] ^ m[31] ^ m[34] ^ m[36] ^ m[38] ^ m[39] ^ m[41] ^ m[43] ^ m[45] ^ m[46] ^ m[49] ^ m[51] ^ m[52] ^ m[54] ^ m[55] ^ m[56];
    assign parity[2] = m[0] ^ m[2] ^ m[4] ^ m[6] ^ m[7] ^ m[9] ^ m[12] ^ m[14] ^ m[16] ^ m[18] ^ m[19] ^ m[22] ^ m[24] ^ m[25] ^ m[28] ^ m[30] ^ m[31] ^ m[34] ^ m[35] ^ m[37] ^ m[40] ^ m[42] ^ m[43] ^ m[45] ^ m[46] ^ m[48] ^ m[50] ^ m[53] ^ m[54] ^ m[55] ^ m[56];
    assign parity[3] = m[0] ^ m[2] ^ m[3] ^ m[5] ^ m[8] ^ m[10] ^ m[12] ^ m[14] ^ m[16] ^ m[18] ^ m[19] ^ m[21] ^ m[23] ^ m[26] ^ m[27] ^ m[30] ^ m[32] ^ m[34] ^ m[36] ^ m[37] ^ m[40] ^ m[41] ^ m[43] ^ m[44] ^ m[47] ^ m[48] ^ m[51] ^ m[52] ^ m[53] ^ m[54] ^ m[56];
    assign parity[4] = m[0] ^ m[1] ^ m[3] ^ m[6] ^ m[7] ^ m[10] ^ m[11] ^ m[14] ^ m[15] ^ m[18] ^ m[20] ^ m[21] ^ m[24] ^ m[25] ^ m[28] ^ m[29] ^ m[32] ^ m[33] ^ m[36] ^ m[38] ^ m[40] ^ m[42] ^ m[43] ^ m[45] ^ m[47] ^ m[48] ^ m[51] ^ m[52] ^ m[53] ^ m[55] ^ m[56];
    assign parity[5] = m[0] ^ m[1] ^ m[3] ^ m[5] ^ m[7] ^ m[9] ^ m[11] ^ m[13] ^ m[15] ^ m[17] ^ m[19] ^ m[22] ^ m[23] ^ m[26] ^ m[27] ^ m[30] ^ m[31] ^ m[34] ^ m[35] ^ m[38] ^ m[39] ^ m[42] ^ m[43] ^ m[45] ^ m[47] ^ m[48] ^ m[51] ^ m[52] ^ m[53] ^ m[54] ^ m[55];
    assign parity[6] = m[0] ^ m[1] ^ m[2] ^ m[5] ^ m[6] ^ m[9] ^ m[10] ^ m[13] ^ m[14] ^ m[17] ^ m[18] ^ m[21] ^ m[22] ^ m[25] ^ m[26] ^ m[29] ^ m[30] ^ m[33] ^ m[34] ^ m[37] ^ m[38] ^ m[41] ^ m[42] ^ m[44] ^ m[46] ^ m[47] ^ m[49] ^ m[50] ^ m[51] ^ m[53] ^ m[55];
  end else if ((CodewordWidth == 128) && (MessageWidth == 120)) begin : gen_128_120
    `BR_ASSERT_STATIC(parity_width_matches_a, ParityWidth == 8)
    assign parity[0] = m[1] ^ m[3] ^ m[5] ^ m[7] ^ m[9] ^ m[10] ^ m[13] ^ m[15] ^ m[17] ^ m[19] ^ m[20] ^ m[23] ^ m[25] ^ m[27] ^ m[28] ^ m[31] ^ m[33] ^ m[34] ^ m[37] ^ m[38] ^ m[40] ^ m[43] ^ m[45] ^ m[47] ^ m[49] ^ m[50] ^ m[53] ^ m[55] ^ m[57] ^ m[58] ^ m[61] ^ m[63] ^ m[64] ^ m[67] ^ m[68] ^ m[70] ^ m[73] ^ m[75] ^ m[77] ^ m[78] ^ m[81] ^ m[83] ^ m[84] ^ m[87] ^ m[88] ^ m[90] ^ m[93] ^ m[95] ^ m[96] ^ m[99] ^ m[100] ^ m[102] ^ m[105] ^ m[106] ^ m[108] ^ m[110] ^ m[113] ^ m[114] ^ m[115] ^ m[116] ^ m[117] ^ m[118] ^ m[119];
    assign parity[1] = m[1] ^ m[3] ^ m[5] ^ m[7] ^ m[8] ^ m[11] ^ m[13] ^ m[15] ^ m[17] ^ m[18] ^ m[21] ^ m[23] ^ m[25] ^ m[26] ^ m[29] ^ m[31] ^ m[32] ^ m[35] ^ m[36] ^ m[39] ^ m[40] ^ m[43] ^ m[45] ^ m[47] ^ m[48] ^ m[51] ^ m[53] ^ m[55] ^ m[56] ^ m[59] ^ m[61] ^ m[62] ^ m[65] ^ m[66] ^ m[69] ^ m[70] ^ m[73] ^ m[75] ^ m[76] ^ m[79] ^ m[81] ^ m[82] ^ m[85] ^ m[86] ^ m[89] ^ m[90] ^ m[93] ^ m[94] ^ m[97] ^ m[98] ^ m[101] ^ m[102] ^ m[104] ^ m[107] ^ m[108] ^ m[110] ^ m[112] ^ m[114] ^ m[115] ^ m[116] ^ m[117] ^ m[118] ^ m[119];
    assign parity[2] = m[1] ^ m[3] ^ m[5] ^ m[6] ^ m[9] ^ m[11] ^ m[13] ^ m[15] ^ m[16] ^ m[19] ^ m[21] ^ m[23] ^ m[24] ^ m[27] ^ m[29] ^ m[30] ^ m[33] ^ m[35] ^ m[36] ^ m[38] ^ m[41] ^ m[43] ^ m[45] ^ m[46] ^ m[49] ^ m[51] ^ m[53] ^ m[54] ^ m[57] ^ m[59] ^ m[60] ^ m[63] ^ m[65] ^ m[66] ^ m[68] ^ m[71] ^ m[73] ^ m[74] ^ m[77] ^ m[79] ^ m[80] ^ m[83] ^ m[85] ^ m[86] ^ m[88] ^ m[91] ^ m[92] ^ m[95] ^ m[97] ^ m[98] ^ m[100] ^ m[103] ^ m[104] ^ m[106] ^ m[109] ^ m[110] ^ m[112] ^ m[113] ^ m[115] ^ m[116] ^ m[117] ^ m[118] ^ m[119];
    assign parity[3] = m[1] ^ m[3] ^ m[4] ^ m[7] ^ m[9] ^ m[11] ^ m[13] ^ m[14] ^ m[17] ^ m[19] ^ m[21] ^ m[22] ^ m[25] ^ m[27] ^ m[29] ^ m[30] ^ m[32] ^ m[34] ^ m[37] ^ m[39] ^ m[41] ^ m[43] ^ m[44] ^ m[47] ^ m[49] ^ m[51] ^ m[52] ^ m[55] ^ m[57] ^ m[59] ^ m[60] ^ m[62] ^ m[64] ^ m[67] ^ m[69] ^ m[71] ^ m[72] ^ m[75] ^ m[77] ^ m[79] ^ m[80] ^ m[82] ^ m[84] ^ m[87] ^ m[89] ^ m[91] ^ m[92] ^ m[94] ^ m[96] ^ m[99] ^ m[101] ^ m[103] ^ m[104] ^ m[106] ^ m[108] ^ m[111] ^ m[112] ^ m[113] ^ m[114] ^ m[116] ^ m[117] ^ m[118] ^ m[119];
    assign parity[4] = m[1] ^ m[2] ^ m[5] ^ m[7] ^ m[9] ^ m[11] ^ m[12] ^ m[15] ^ m[17] ^ m[19] ^ m[21] ^ m[22] ^ m[24] ^ m[26] ^ m[28] ^ m[31] ^ m[33] ^ m[35] ^ m[37] ^ m[39] ^ m[41] ^ m[42] ^ m[45] ^ m[47] ^ m[49] ^ m[51] ^ m[52] ^ m[54] ^ m[56] ^ m[58] ^ m[61] ^ m[63] ^ m[65] ^ m[67] ^ m[69] ^ m[71] ^ m[72] ^ m[74] ^ m[76] ^ m[78] ^ m[81] ^ m[83] ^ m[85] ^ m[87] ^ m[89] ^ m[91] ^ m[92] ^ m[94] ^ m[96] ^ m[98] ^ m[100] ^ m[102] ^ m[105] ^ m[107] ^ m[109] ^ m[111] ^ m[112] ^ m[113] ^ m[114] ^ m[115] ^ m[117] ^ m[118] ^ m[119];
    assign parity[5] = m[0] ^ m[3] ^ m[5] ^ m[7] ^ m[9] ^ m[11] ^ m[12] ^ m[14] ^ m[16] ^ m[18] ^ m[20] ^ m[23] ^ m[25] ^ m[27] ^ m[29] ^ m[31] ^ m[33] ^ m[35] ^ m[37] ^ m[39] ^ m[41] ^ m[42] ^ m[44] ^ m[46] ^ m[48] ^ m[50] ^ m[53] ^ m[55] ^ m[57] ^ m[59] ^ m[61] ^ m[63] ^ m[65] ^ m[67] ^ m[69] ^ m[71] ^ m[72] ^ m[74] ^ m[76] ^ m[78] ^ m[80] ^ m[82] ^ m[84] ^ m[86] ^ m[88] ^ m[90] ^ m[93] ^ m[95] ^ m[97] ^ m[99] ^ m[101] ^ m[103] ^ m[105] ^ m[107] ^ m[109] ^ m[111] ^ m[112] ^ m[113] ^ m[114] ^ m[115] ^ m[116] ^ m[118] ^ m[119];
    assign parity[6] = m[0] ^ m[2] ^ m[4] ^ m[6] ^ m[8] ^ m[10] ^ m[13] ^ m[15] ^ m[17] ^ m[19] ^ m[21] ^ m[23] ^ m[25] ^ m[27] ^ m[29] ^ m[31] ^ m[33] ^ m[35] ^ m[37] ^ m[39] ^ m[41] ^ m[42] ^ m[44] ^ m[46] ^ m[48] ^ m[50] ^ m[52] ^ m[54] ^ m[56] ^ m[58] ^ m[60] ^ m[62] ^ m[64] ^ m[66] ^ m[68] ^ m[70] ^ m[73] ^ m[75] ^ m[77] ^ m[79] ^ m[81] ^ m[83] ^ m[85] ^ m[87] ^ m[89] ^ m[91] ^ m[93] ^ m[95] ^ m[97] ^ m[99] ^ m[101] ^ m[103] ^ m[105] ^ m[107] ^ m[109] ^ m[111] ^ m[112] ^ m[113] ^ m[114] ^ m[115] ^ m[116] ^ m[117] ^ m[119];
    assign parity[7] = m[0] ^ m[2] ^ m[4] ^ m[6] ^ m[8] ^ m[10] ^ m[12] ^ m[14] ^ m[16] ^ m[18] ^ m[20] ^ m[22] ^ m[24] ^ m[26] ^ m[28] ^ m[30] ^ m[32] ^ m[34] ^ m[36] ^ m[38] ^ m[40] ^ m[43] ^ m[45] ^ m[47] ^ m[49] ^ m[51] ^ m[53] ^ m[55] ^ m[57] ^ m[59] ^ m[61] ^ m[63] ^ m[65] ^ m[67] ^ m[69] ^ m[71] ^ m[73] ^ m[75] ^ m[77] ^ m[79] ^ m[81] ^ m[83] ^ m[85] ^ m[87] ^ m[89] ^ m[91] ^ m[93] ^ m[95] ^ m[97] ^ m[99] ^ m[101] ^ m[103] ^ m[105] ^ m[107] ^ m[109] ^ m[111] ^ m[112] ^ m[113] ^ m[114] ^ m[115] ^ m[116] ^ m[117] ^ m[118];
  end else if ((CodewordWidth == 256) && (MessageWidth == 247)) begin : gen_256_247
    `BR_ASSERT_STATIC(parity_width_matches_a, ParityWidth == 9)
    assign parity[0] = m[0] ^ m[2] ^ m[4] ^ m[6] ^ m[8] ^ m[10] ^ m[12] ^ m[14] ^ m[16] ^ m[18] ^ m[20] ^ m[22] ^ m[23] ^ m[25] ^ m[28] ^ m[30] ^ m[32] ^ m[34] ^ m[36] ^ m[38] ^ m[40] ^ m[42] ^ m[43] ^ m[46] ^ m[48] ^ m[49] ^ m[52] ^ m[54] ^ m[56] ^ m[58] ^ m[59] ^ m[62] ^ m[64] ^ m[66] ^ m[68] ^ m[69] ^ m[71] ^ m[74] ^ m[76] ^ m[78] ^ m[79] ^ m[82] ^ m[83] ^ m[85] ^ m[88] ^ m[90] ^ m[92] ^ m[94] ^ m[96] ^ m[97] ^ m[100] ^ m[102] ^ m[103] ^ m[105] ^ m[108] ^ m[109] ^ m[112] ^ m[115] ^ m[117] ^ m[119] ^ m[120] ^ m[124] ^ m[126] ^ m[129] ^ m[130] ^ m[132] ^ m[135] ^ m[137] ^ m[139] ^ m[143] ^ m[144] ^ m[147] ^ m[148] ^ m[152] ^ m[153] ^ m[155] ^ m[158] ^ m[159] ^ m[161] ^ m[162] ^ m[166] ^ m[168] ^ m[170] ^ m[171] ^ m[173] ^ m[175] ^ m[177] ^ m[178] ^ m[180] ^ m[181] ^ m[183] ^ m[185] ^ m[187] ^ m[188] ^ m[190] ^ m[193] ^ m[194] ^ m[195] ^ m[198] ^ m[200] ^ m[201] ^ m[203] ^ m[205] ^ m[206] ^ m[209] ^ m[211] ^ m[212] ^ m[214] ^ m[215] ^ m[218] ^ m[220] ^ m[221] ^ m[223] ^ m[225] ^ m[227] ^ m[228] ^ m[230] ^ m[232] ^ m[234] ^ m[236] ^ m[237] ^ m[239] ^ m[240] ^ m[242] ^ m[243] ^ m[245] ^ m[246];
    assign parity[1] = m[0] ^ m[2] ^ m[4] ^ m[6] ^ m[8] ^ m[10] ^ m[12] ^ m[14] ^ m[16] ^ m[18] ^ m[19] ^ m[21] ^ m[24] ^ m[26] ^ m[28] ^ m[30] ^ m[32] ^ m[34] ^ m[36] ^ m[38] ^ m[39] ^ m[42] ^ m[44] ^ m[45] ^ m[48] ^ m[50] ^ m[52] ^ m[54] ^ m[55] ^ m[58] ^ m[60] ^ m[62] ^ m[64] ^ m[65] ^ m[67] ^ m[70] ^ m[72] ^ m[74] ^ m[75] ^ m[78] ^ m[80] ^ m[81] ^ m[83] ^ m[86] ^ m[88] ^ m[90] ^ m[92] ^ m[93] ^ m[96] ^ m[98] ^ m[99] ^ m[101] ^ m[104] ^ m[106] ^ m[108] ^ m[109] ^ m[112] ^ m[113] ^ m[117] ^ m[119] ^ m[121] ^ m[123] ^ m[126] ^ m[128] ^ m[131] ^ m[133] ^ m[134] ^ m[138] ^ m[140] ^ m[141] ^ m[144] ^ m[146] ^ m[148] ^ m[150] ^ m[153] ^ m[154] ^ m[156] ^ m[159] ^ m[161] ^ m[163] ^ m[164] ^ m[168] ^ m[170] ^ m[171] ^ m[173] ^ m[175] ^ m[177] ^ m[178] ^ m[179] ^ m[181] ^ m[182] ^ m[184] ^ m[186] ^ m[189] ^ m[191] ^ m[193] ^ m[194] ^ m[196] ^ m[198] ^ m[199] ^ m[201] ^ m[202] ^ m[204] ^ m[207] ^ m[208] ^ m[210] ^ m[212] ^ m[214] ^ m[216] ^ m[218] ^ m[219] ^ m[222] ^ m[224] ^ m[226] ^ m[227] ^ m[229] ^ m[230] ^ m[233] ^ m[234] ^ m[236] ^ m[238] ^ m[239] ^ m[241] ^ m[242] ^ m[244] ^ m[245] ^ m[246];
    assign parity[2] = m[0] ^ m[2] ^ m[4] ^ m[6] ^ m[8] ^ m[10] ^ m[12] ^ m[14] ^ m[15] ^ m[17] ^ m[20] ^ m[22] ^ m[24] ^ m[26] ^ m[28] ^ m[30] ^ m[32] ^ m[34] ^ m[35] ^ m[38] ^ m[40] ^ m[41] ^ m[44] ^ m[46] ^ m[48] ^ m[50] ^ m[51] ^ m[54] ^ m[56] ^ m[58] ^ m[60] ^ m[61] ^ m[63] ^ m[66] ^ m[68] ^ m[70] ^ m[72] ^ m[74] ^ m[75] ^ m[77] ^ m[79] ^ m[82] ^ m[84] ^ m[86] ^ m[88] ^ m[89] ^ m[92] ^ m[94] ^ m[95] ^ m[98] ^ m[100] ^ m[101] ^ m[104] ^ m[105] ^ m[108] ^ m[110] ^ m[111] ^ m[114] ^ m[116] ^ m[119] ^ m[122] ^ m[124] ^ m[125] ^ m[127] ^ m[131] ^ m[133] ^ m[135] ^ m[138] ^ m[140] ^ m[141] ^ m[143] ^ m[146] ^ m[149] ^ m[150] ^ m[152] ^ m[154] ^ m[157] ^ m[158] ^ m[161] ^ m[162] ^ m[165] ^ m[167] ^ m[170] ^ m[171] ^ m[172] ^ m[174] ^ m[176] ^ m[178] ^ m[180] ^ m[181] ^ m[183] ^ m[185] ^ m[187] ^ m[189] ^ m[191] ^ m[192] ^ m[194] ^ m[196] ^ m[197] ^ m[200] ^ m[201] ^ m[203] ^ m[204] ^ m[207] ^ m[208] ^ m[211] ^ m[212] ^ m[213] ^ m[215] ^ m[217] ^ m[220] ^ m[222] ^ m[223] ^ m[225] ^ m[226] ^ m[229] ^ m[231] ^ m[232] ^ m[234] ^ m[235] ^ m[238] ^ m[239] ^ m[240] ^ m[241] ^ m[243] ^ m[244] ^ m[245];
    assign parity[3] = m[0] ^ m[2] ^ m[4] ^ m[6] ^ m[8] ^ m[10] ^ m[11] ^ m[13] ^ m[16] ^ m[18] ^ m[20] ^ m[22] ^ m[24] ^ m[26] ^ m[28] ^ m[30] ^ m[31] ^ m[34] ^ m[36] ^ m[37] ^ m[40] ^ m[42] ^ m[44] ^ m[46] ^ m[47] ^ m[50] ^ m[52] ^ m[54] ^ m[56] ^ m[57] ^ m[60] ^ m[62] ^ m[63] ^ m[66] ^ m[67] ^ m[70] ^ m[71] ^ m[73] ^ m[76] ^ m[78] ^ m[80] ^ m[82] ^ m[84] ^ m[86] ^ m[88] ^ m[89] ^ m[91] ^ m[93] ^ m[96] ^ m[97] ^ m[100] ^ m[102] ^ m[104] ^ m[106] ^ m[107] ^ m[110] ^ m[112] ^ m[114] ^ m[116] ^ m[118] ^ m[121] ^ m[123] ^ m[126] ^ m[127] ^ m[130] ^ m[133] ^ m[134] ^ m[137] ^ m[139] ^ m[142] ^ m[145] ^ m[147] ^ m[150] ^ m[151] ^ m[155] ^ m[157] ^ m[158] ^ m[159] ^ m[160] ^ m[162] ^ m[166] ^ m[168] ^ m[169] ^ m[171] ^ m[172] ^ m[175] ^ m[176] ^ m[178] ^ m[180] ^ m[181] ^ m[182] ^ m[185] ^ m[186] ^ m[189] ^ m[191] ^ m[192] ^ m[194] ^ m[196] ^ m[197] ^ m[199] ^ m[201] ^ m[202] ^ m[205] ^ m[206] ^ m[209] ^ m[210] ^ m[211] ^ m[213] ^ m[216] ^ m[217] ^ m[219] ^ m[221] ^ m[224] ^ m[226] ^ m[227] ^ m[228] ^ m[231] ^ m[232] ^ m[233] ^ m[235] ^ m[237] ^ m[238] ^ m[240] ^ m[242] ^ m[243] ^ m[244] ^ m[246];
    assign parity[4] = m[0] ^ m[2] ^ m[4] ^ m[6] ^ m[7] ^ m[9] ^ m[12] ^ m[14] ^ m[16] ^ m[18] ^ m[20] ^ m[22] ^ m[24] ^ m[26] ^ m[27] ^ m[30] ^ m[32] ^ m[33] ^ m[36] ^ m[38] ^ m[40] ^ m[42] ^ m[44] ^ m[46] ^ m[47] ^ m[50] ^ m[51] ^ m[53] ^ m[55] ^ m[58] ^ m[59] ^ m[62] ^ m[64] ^ m[66] ^ m[68] ^ m[70] ^ m[72] ^ m[73] ^ m[76] ^ m[77] ^ m[80] ^ m[81] ^ m[84] ^ m[85] ^ m[87] ^ m[90] ^ m[92] ^ m[94] ^ m[96] ^ m[98] ^ m[100] ^ m[102] ^ m[104] ^ m[106] ^ m[107] ^ m[110] ^ m[111] ^ m[113] ^ m[116] ^ m[118] ^ m[120] ^ m[123] ^ m[125] ^ m[128] ^ m[129] ^ m[132] ^ m[136] ^ m[137] ^ m[140] ^ m[142] ^ m[145] ^ m[147] ^ m[149] ^ m[152] ^ m[153] ^ m[154] ^ m[158] ^ m[160] ^ m[163] ^ m[164] ^ m[165] ^ m[167] ^ m[169] ^ m[171] ^ m[173] ^ m[174] ^ m[176] ^ m[178] ^ m[179] ^ m[181] ^ m[183] ^ m[184] ^ m[186] ^ m[188] ^ m[190] ^ m[192] ^ m[193] ^ m[195] ^ m[196] ^ m[199] ^ m[200] ^ m[203] ^ m[205] ^ m[206] ^ m[208] ^ m[211] ^ m[212] ^ m[213] ^ m[214] ^ m[216] ^ m[220] ^ m[222] ^ m[224] ^ m[225] ^ m[227] ^ m[228] ^ m[229] ^ m[230] ^ m[231] ^ m[233] ^ m[235] ^ m[236] ^ m[237] ^ m[241] ^ m[244] ^ m[245] ^ m[246];
    assign parity[5] = m[0] ^ m[2] ^ m[3] ^ m[5] ^ m[8] ^ m[10] ^ m[12] ^ m[14] ^ m[16] ^ m[18] ^ m[20] ^ m[22] ^ m[24] ^ m[26] ^ m[27] ^ m[29] ^ m[31] ^ m[34] ^ m[35] ^ m[38] ^ m[39] ^ m[42] ^ m[43] ^ m[46] ^ m[48] ^ m[50] ^ m[52] ^ m[53] ^ m[56] ^ m[57] ^ m[60] ^ m[61] ^ m[64] ^ m[65] ^ m[68] ^ m[69] ^ m[72] ^ m[74] ^ m[76] ^ m[78] ^ m[80] ^ m[82] ^ m[84] ^ m[86] ^ m[87] ^ m[90] ^ m[91] ^ m[94] ^ m[95] ^ m[98] ^ m[99] ^ m[102] ^ m[103] ^ m[106] ^ m[108] ^ m[110] ^ m[112] ^ m[114] ^ m[115] ^ m[118] ^ m[121] ^ m[122] ^ m[125] ^ m[128] ^ m[130] ^ m[132] ^ m[135] ^ m[136] ^ m[138] ^ m[142] ^ m[144] ^ m[146] ^ m[149] ^ m[151] ^ m[156] ^ m[157] ^ m[158] ^ m[160] ^ m[164] ^ m[165] ^ m[166] ^ m[168] ^ m[169] ^ m[171] ^ m[173] ^ m[174] ^ m[176] ^ m[177] ^ m[179] ^ m[181] ^ m[183] ^ m[184] ^ m[186] ^ m[187] ^ m[188] ^ m[190] ^ m[191] ^ m[194] ^ m[195] ^ m[197] ^ m[198] ^ m[202] ^ m[204] ^ m[206] ^ m[207] ^ m[208] ^ m[209] ^ m[210] ^ m[212] ^ m[215] ^ m[217] ^ m[218] ^ m[219] ^ m[221] ^ m[223] ^ m[225] ^ m[226] ^ m[230] ^ m[232] ^ m[233] ^ m[235] ^ m[237] ^ m[239] ^ m[241] ^ m[243] ^ m[244] ^ m[246];
    assign parity[6] = m[0] ^ m[1] ^ m[3] ^ m[6] ^ m[7] ^ m[10] ^ m[11] ^ m[14] ^ m[15] ^ m[18] ^ m[19] ^ m[22] ^ m[23] ^ m[26] ^ m[28] ^ m[29] ^ m[32] ^ m[33] ^ m[36] ^ m[37] ^ m[40] ^ m[41] ^ m[44] ^ m[45] ^ m[48] ^ m[49] ^ m[52] ^ m[54] ^ m[56] ^ m[58] ^ m[60] ^ m[62] ^ m[64] ^ m[66] ^ m[68] ^ m[70] ^ m[72] ^ m[74] ^ m[76] ^ m[78] ^ m[80] ^ m[82] ^ m[84] ^ m[86] ^ m[87] ^ m[90] ^ m[91] ^ m[94] ^ m[95] ^ m[98] ^ m[99] ^ m[102] ^ m[103] ^ m[106] ^ m[107] ^ m[110] ^ m[111] ^ m[113] ^ m[115] ^ m[117] ^ m[120] ^ m[122] ^ m[124] ^ m[127] ^ m[129] ^ m[131] ^ m[134] ^ m[136] ^ m[139] ^ m[141] ^ m[143] ^ m[145] ^ m[148] ^ m[151] ^ m[155] ^ m[156] ^ m[158] ^ m[160] ^ m[163] ^ m[165] ^ m[166] ^ m[167] ^ m[169] ^ m[170] ^ m[172] ^ m[174] ^ m[175] ^ m[178] ^ m[179] ^ m[181] ^ m[182] ^ m[184] ^ m[185] ^ m[189] ^ m[190] ^ m[192] ^ m[194] ^ m[195] ^ m[197] ^ m[198] ^ m[199] ^ m[202] ^ m[203] ^ m[204] ^ m[205] ^ m[207] ^ m[212] ^ m[214] ^ m[215] ^ m[217] ^ m[218] ^ m[219] ^ m[220] ^ m[221] ^ m[222] ^ m[223] ^ m[224] ^ m[228] ^ m[229] ^ m[231] ^ m[234] ^ m[236] ^ m[238] ^ m[240] ^ m[242] ^ m[244] ^ m[246];
    assign parity[7] = m[0] ^ m[1] ^ m[3] ^ m[5] ^ m[7] ^ m[9] ^ m[11] ^ m[13] ^ m[15] ^ m[17] ^ m[19] ^ m[21] ^ m[23] ^ m[25] ^ m[27] ^ m[30] ^ m[31] ^ m[34] ^ m[35] ^ m[38] ^ m[39] ^ m[42] ^ m[43] ^ m[46] ^ m[47] ^ m[50] ^ m[51] ^ m[54] ^ m[55] ^ m[58] ^ m[59] ^ m[62] ^ m[63] ^ m[66] ^ m[67] ^ m[70] ^ m[71] ^ m[74] ^ m[75] ^ m[78] ^ m[79] ^ m[82] ^ m[83] ^ m[86] ^ m[88] ^ m[90] ^ m[92] ^ m[94] ^ m[96] ^ m[98] ^ m[100] ^ m[102] ^ m[104] ^ m[106] ^ m[108] ^ m[110] ^ m[112] ^ m[115] ^ m[117] ^ m[119] ^ m[122] ^ m[124] ^ m[126] ^ m[129] ^ m[131] ^ m[133] ^ m[136] ^ m[138] ^ m[140] ^ m[142] ^ m[145] ^ m[147] ^ m[149] ^ m[151] ^ m[155] ^ m[156] ^ m[157] ^ m[158] ^ m[163] ^ m[164] ^ m[166] ^ m[167] ^ m[169] ^ m[171] ^ m[172] ^ m[174] ^ m[176] ^ m[177] ^ m[178] ^ m[180] ^ m[182] ^ m[184] ^ m[186] ^ m[187] ^ m[188] ^ m[190] ^ m[192] ^ m[193] ^ m[194] ^ m[197] ^ m[199] ^ m[200] ^ m[202] ^ m[204] ^ m[206] ^ m[208] ^ m[209] ^ m[210] ^ m[212] ^ m[213] ^ m[215] ^ m[216] ^ m[218] ^ m[220] ^ m[222] ^ m[225] ^ m[226] ^ m[228] ^ m[230] ^ m[232] ^ m[234] ^ m[236] ^ m[238] ^ m[240] ^ m[242] ^ m[244] ^ m[246];
    assign parity[8] = m[0] ^ m[1] ^ m[2] ^ m[5] ^ m[6] ^ m[9] ^ m[10] ^ m[13] ^ m[14] ^ m[17] ^ m[18] ^ m[21] ^ m[22] ^ m[25] ^ m[26] ^ m[29] ^ m[30] ^ m[33] ^ m[34] ^ m[37] ^ m[38] ^ m[41] ^ m[42] ^ m[45] ^ m[46] ^ m[49] ^ m[50] ^ m[53] ^ m[54] ^ m[57] ^ m[58] ^ m[61] ^ m[62] ^ m[65] ^ m[66] ^ m[69] ^ m[70] ^ m[73] ^ m[74] ^ m[77] ^ m[78] ^ m[81] ^ m[82] ^ m[85] ^ m[86] ^ m[89] ^ m[90] ^ m[93] ^ m[94] ^ m[97] ^ m[98] ^ m[101] ^ m[102] ^ m[105] ^ m[106] ^ m[109] ^ m[110] ^ m[115] ^ m[117] ^ m[119] ^ m[122] ^ m[124] ^ m[126] ^ m[129] ^ m[131] ^ m[133] ^ m[136] ^ m[138] ^ m[140] ^ m[142] ^ m[145] ^ m[147] ^ m[149] ^ m[151] ^ m[155] ^ m[156] ^ m[157] ^ m[160] ^ m[163] ^ m[164] ^ m[165] ^ m[167] ^ m[168] ^ m[170] ^ m[172] ^ m[173] ^ m[175] ^ m[177] ^ m[179] ^ m[180] ^ m[182] ^ m[183] ^ m[185] ^ m[187] ^ m[188] ^ m[189] ^ m[191] ^ m[193] ^ m[195] ^ m[196] ^ m[198] ^ m[200] ^ m[201] ^ m[203] ^ m[205] ^ m[207] ^ m[209] ^ m[210] ^ m[211] ^ m[213] ^ m[214] ^ m[216] ^ m[217] ^ m[219] ^ m[221] ^ m[223] ^ m[224] ^ m[227] ^ m[229] ^ m[231] ^ m[233] ^ m[235] ^ m[237] ^ m[239] ^ m[241] ^ m[243] ^ m[245];
  end else if ((CodewordWidth == 512) && (MessageWidth == 502)) begin : gen_512_502
    `BR_ASSERT_STATIC(parity_width_matches_a, ParityWidth == 10)
    assign parity[0] = m[1] ^ m[3] ^ m[5] ^ m[7] ^ m[9] ^ m[11] ^ m[13] ^ m[14] ^ m[17] ^ m[19] ^ m[21] ^ m[23] ^ m[25] ^ m[27] ^ m[28] ^ m[31] ^ m[33] ^ m[35] ^ m[37] ^ m[39] ^ m[40] ^ m[43] ^ m[45] ^ m[47] ^ m[49] ^ m[50] ^ m[53] ^ m[55] ^ m[57] ^ m[58] ^ m[61] ^ m[63] ^ m[64] ^ m[67] ^ m[68] ^ m[70] ^ m[73] ^ m[75] ^ m[77] ^ m[79] ^ m[81] ^ m[83] ^ m[84] ^ m[87] ^ m[89] ^ m[91] ^ m[93] ^ m[95] ^ m[96] ^ m[99] ^ m[101] ^ m[103] ^ m[105] ^ m[106] ^ m[109] ^ m[111] ^ m[113] ^ m[114] ^ m[117] ^ m[119] ^ m[120] ^ m[123] ^ m[124] ^ m[126] ^ m[129] ^ m[131] ^ m[133] ^ m[135] ^ m[137] ^ m[138] ^ m[141] ^ m[143] ^ m[145] ^ m[147] ^ m[148] ^ m[151] ^ m[153] ^ m[155] ^ m[156] ^ m[159] ^ m[161] ^ m[162] ^ m[165] ^ m[166] ^ m[168] ^ m[171] ^ m[173] ^ m[175] ^ m[177] ^ m[178] ^ m[181] ^ m[183] ^ m[185] ^ m[186] ^ m[189] ^ m[191] ^ m[192] ^ m[195] ^ m[196] ^ m[198] ^ m[201] ^ m[203] ^ m[205] ^ m[206] ^ m[209] ^ m[211] ^ m[212] ^ m[215] ^ m[216] ^ m[218] ^ m[221] ^ m[223] ^ m[224] ^ m[227] ^ m[228] ^ m[230] ^ m[233] ^ m[234] ^ m[236] ^ m[238] ^ m[241] ^ m[243] ^ m[245] ^ m[247] ^ m[249] ^ m[250] ^ m[253] ^ m[255] ^ m[257] ^ m[259] ^ m[260] ^ m[263] ^ m[265] ^ m[267] ^ m[268] ^ m[271] ^ m[273] ^ m[274] ^ m[277] ^ m[278] ^ m[280] ^ m[283] ^ m[285] ^ m[287] ^ m[289] ^ m[290] ^ m[293] ^ m[295] ^ m[297] ^ m[298] ^ m[301] ^ m[303] ^ m[304] ^ m[307] ^ m[308] ^ m[310] ^ m[313] ^ m[315] ^ m[317] ^ m[318] ^ m[321] ^ m[323] ^ m[324] ^ m[327] ^ m[328] ^ m[330] ^ m[333] ^ m[335] ^ m[336] ^ m[339] ^ m[340] ^ m[342] ^ m[345] ^ m[346] ^ m[348] ^ m[350] ^ m[353] ^ m[355] ^ m[357] ^ m[359] ^ m[360] ^ m[363] ^ m[365] ^ m[367] ^ m[368] ^ m[371] ^ m[373] ^ m[374] ^ m[377] ^ m[378] ^ m[380] ^ m[383] ^ m[385] ^ m[387] ^ m[388] ^ m[391] ^ m[393] ^ m[394] ^ m[397] ^ m[398] ^ m[400] ^ m[403] ^ m[405] ^ m[406] ^ m[409] ^ m[410] ^ m[412] ^ m[415] ^ m[416] ^ m[418] ^ m[420] ^ m[423] ^ m[425] ^ m[427] ^ m[428] ^ m[431] ^ m[433] ^ m[434] ^ m[437] ^ m[438] ^ m[440] ^ m[443] ^ m[445] ^ m[446] ^ m[449] ^ m[450] ^ m[452] ^ m[455] ^ m[456] ^ m[458] ^ m[460] ^ m[463] ^ m[465] ^ m[466] ^ m[469] ^ m[470] ^ m[472] ^ m[475] ^ m[476] ^ m[478] ^ m[480] ^ m[483] ^ m[484] ^ m[486] ^ m[488] ^ m[490] ^ m[493] ^ m[494] ^ m[495] ^ m[496] ^ m[497] ^ m[498] ^ m[499] ^ m[500] ^ m[501];
    assign parity[1] = m[1] ^ m[3] ^ m[5] ^ m[7] ^ m[9] ^ m[11] ^ m[12] ^ m[15] ^ m[17] ^ m[19] ^ m[21] ^ m[23] ^ m[25] ^ m[26] ^ m[29] ^ m[31] ^ m[33] ^ m[35] ^ m[37] ^ m[38] ^ m[41] ^ m[43] ^ m[45] ^ m[47] ^ m[48] ^ m[51] ^ m[53] ^ m[55] ^ m[56] ^ m[59] ^ m[61] ^ m[62] ^ m[65] ^ m[66] ^ m[69] ^ m[70] ^ m[73] ^ m[75] ^ m[77] ^ m[79] ^ m[81] ^ m[82] ^ m[85] ^ m[87] ^ m[89] ^ m[91] ^ m[93] ^ m[94] ^ m[97] ^ m[99] ^ m[101] ^ m[103] ^ m[104] ^ m[107] ^ m[109] ^ m[111] ^ m[112] ^ m[115] ^ m[117] ^ m[118] ^ m[121] ^ m[122] ^ m[125] ^ m[126] ^ m[129] ^ m[131] ^ m[133] ^ m[135] ^ m[136] ^ m[139] ^ m[141] ^ m[143] ^ m[145] ^ m[146] ^ m[149] ^ m[151] ^ m[153] ^ m[154] ^ m[157] ^ m[159] ^ m[160] ^ m[163] ^ m[164] ^ m[167] ^ m[168] ^ m[171] ^ m[173] ^ m[175] ^ m[176] ^ m[179] ^ m[181] ^ m[183] ^ m[184] ^ m[187] ^ m[189] ^ m[190] ^ m[193] ^ m[194] ^ m[197] ^ m[198] ^ m[201] ^ m[203] ^ m[204] ^ m[207] ^ m[209] ^ m[210] ^ m[213] ^ m[214] ^ m[217] ^ m[218] ^ m[221] ^ m[222] ^ m[225] ^ m[226] ^ m[229] ^ m[230] ^ m[232] ^ m[235] ^ m[236] ^ m[238] ^ m[241] ^ m[243] ^ m[245] ^ m[247] ^ m[248] ^ m[251] ^ m[253] ^ m[255] ^ m[257] ^ m[258] ^ m[261] ^ m[263] ^ m[265] ^ m[266] ^ m[269] ^ m[271] ^ m[272] ^ m[275] ^ m[276] ^ m[279] ^ m[280] ^ m[283] ^ m[285] ^ m[287] ^ m[288] ^ m[291] ^ m[293] ^ m[295] ^ m[296] ^ m[299] ^ m[301] ^ m[302] ^ m[305] ^ m[306] ^ m[309] ^ m[310] ^ m[313] ^ m[315] ^ m[316] ^ m[319] ^ m[321] ^ m[322] ^ m[325] ^ m[326] ^ m[329] ^ m[330] ^ m[333] ^ m[334] ^ m[337] ^ m[338] ^ m[341] ^ m[342] ^ m[344] ^ m[347] ^ m[348] ^ m[350] ^ m[353] ^ m[355] ^ m[357] ^ m[358] ^ m[361] ^ m[363] ^ m[365] ^ m[366] ^ m[369] ^ m[371] ^ m[372] ^ m[375] ^ m[376] ^ m[379] ^ m[380] ^ m[383] ^ m[385] ^ m[386] ^ m[389] ^ m[391] ^ m[392] ^ m[395] ^ m[396] ^ m[399] ^ m[400] ^ m[403] ^ m[404] ^ m[407] ^ m[408] ^ m[411] ^ m[412] ^ m[414] ^ m[417] ^ m[418] ^ m[420] ^ m[423] ^ m[425] ^ m[426] ^ m[429] ^ m[431] ^ m[432] ^ m[435] ^ m[436] ^ m[439] ^ m[440] ^ m[443] ^ m[444] ^ m[447] ^ m[448] ^ m[451] ^ m[452] ^ m[454] ^ m[457] ^ m[458] ^ m[460] ^ m[463] ^ m[464] ^ m[467] ^ m[468] ^ m[471] ^ m[472] ^ m[474] ^ m[477] ^ m[478] ^ m[480] ^ m[482] ^ m[485] ^ m[486] ^ m[488] ^ m[490] ^ m[492] ^ m[494] ^ m[495] ^ m[496] ^ m[497] ^ m[498] ^ m[499] ^ m[500] ^ m[501];
    assign parity[2] = m[1] ^ m[3] ^ m[5] ^ m[7] ^ m[9] ^ m[10] ^ m[13] ^ m[15] ^ m[17] ^ m[19] ^ m[21] ^ m[23] ^ m[24] ^ m[27] ^ m[29] ^ m[31] ^ m[33] ^ m[35] ^ m[36] ^ m[39] ^ m[41] ^ m[43] ^ m[45] ^ m[46] ^ m[49] ^ m[51] ^ m[53] ^ m[54] ^ m[57] ^ m[59] ^ m[60] ^ m[63] ^ m[65] ^ m[66] ^ m[68] ^ m[71] ^ m[73] ^ m[75] ^ m[77] ^ m[79] ^ m[80] ^ m[83] ^ m[85] ^ m[87] ^ m[89] ^ m[91] ^ m[92] ^ m[95] ^ m[97] ^ m[99] ^ m[101] ^ m[102] ^ m[105] ^ m[107] ^ m[109] ^ m[110] ^ m[113] ^ m[115] ^ m[116] ^ m[119] ^ m[121] ^ m[122] ^ m[124] ^ m[127] ^ m[129] ^ m[131] ^ m[133] ^ m[134] ^ m[137] ^ m[139] ^ m[141] ^ m[143] ^ m[144] ^ m[147] ^ m[149] ^ m[151] ^ m[152] ^ m[155] ^ m[157] ^ m[158] ^ m[161] ^ m[163] ^ m[164] ^ m[166] ^ m[169] ^ m[171] ^ m[173] ^ m[174] ^ m[177] ^ m[179] ^ m[181] ^ m[182] ^ m[185] ^ m[187] ^ m[188] ^ m[191] ^ m[193] ^ m[194] ^ m[196] ^ m[199] ^ m[201] ^ m[202] ^ m[205] ^ m[207] ^ m[208] ^ m[211] ^ m[213] ^ m[214] ^ m[216] ^ m[219] ^ m[220] ^ m[223] ^ m[225] ^ m[226] ^ m[228] ^ m[231] ^ m[232] ^ m[234] ^ m[237] ^ m[238] ^ m[241] ^ m[243] ^ m[245] ^ m[246] ^ m[249] ^ m[251] ^ m[253] ^ m[255] ^ m[256] ^ m[259] ^ m[261] ^ m[263] ^ m[264] ^ m[267] ^ m[269] ^ m[270] ^ m[273] ^ m[275] ^ m[276] ^ m[278] ^ m[281] ^ m[283] ^ m[285] ^ m[286] ^ m[289] ^ m[291] ^ m[293] ^ m[294] ^ m[297] ^ m[299] ^ m[300] ^ m[303] ^ m[305] ^ m[306] ^ m[308] ^ m[311] ^ m[313] ^ m[314] ^ m[317] ^ m[319] ^ m[320] ^ m[323] ^ m[325] ^ m[326] ^ m[328] ^ m[331] ^ m[332] ^ m[335] ^ m[337] ^ m[338] ^ m[340] ^ m[343] ^ m[344] ^ m[346] ^ m[349] ^ m[350] ^ m[353] ^ m[355] ^ m[356] ^ m[359] ^ m[361] ^ m[363] ^ m[364] ^ m[367] ^ m[369] ^ m[370] ^ m[373] ^ m[375] ^ m[376] ^ m[378] ^ m[381] ^ m[383] ^ m[384] ^ m[387] ^ m[389] ^ m[390] ^ m[393] ^ m[395] ^ m[396] ^ m[398] ^ m[401] ^ m[402] ^ m[405] ^ m[407] ^ m[408] ^ m[410] ^ m[413] ^ m[414] ^ m[416] ^ m[419] ^ m[420] ^ m[423] ^ m[424] ^ m[427] ^ m[429] ^ m[430] ^ m[433] ^ m[435] ^ m[436] ^ m[438] ^ m[441] ^ m[442] ^ m[445] ^ m[447] ^ m[448] ^ m[450] ^ m[453] ^ m[454] ^ m[456] ^ m[459] ^ m[460] ^ m[462] ^ m[465] ^ m[467] ^ m[468] ^ m[470] ^ m[473] ^ m[474] ^ m[476] ^ m[479] ^ m[480] ^ m[482] ^ m[484] ^ m[487] ^ m[488] ^ m[490] ^ m[492] ^ m[493] ^ m[495] ^ m[496] ^ m[497] ^ m[498] ^ m[499] ^ m[500] ^ m[501];
    assign parity[3] = m[1] ^ m[3] ^ m[5] ^ m[7] ^ m[8] ^ m[11] ^ m[13] ^ m[15] ^ m[17] ^ m[19] ^ m[21] ^ m[22] ^ m[25] ^ m[27] ^ m[29] ^ m[31] ^ m[33] ^ m[34] ^ m[37] ^ m[39] ^ m[41] ^ m[43] ^ m[44] ^ m[47] ^ m[49] ^ m[51] ^ m[52] ^ m[55] ^ m[57] ^ m[59] ^ m[60] ^ m[62] ^ m[64] ^ m[67] ^ m[69] ^ m[71] ^ m[73] ^ m[75] ^ m[77] ^ m[78] ^ m[81] ^ m[83] ^ m[85] ^ m[87] ^ m[89] ^ m[90] ^ m[93] ^ m[95] ^ m[97] ^ m[99] ^ m[100] ^ m[103] ^ m[105] ^ m[107] ^ m[108] ^ m[111] ^ m[113] ^ m[115] ^ m[116] ^ m[118] ^ m[120] ^ m[123] ^ m[125] ^ m[127] ^ m[129] ^ m[131] ^ m[132] ^ m[135] ^ m[137] ^ m[139] ^ m[141] ^ m[142] ^ m[145] ^ m[147] ^ m[149] ^ m[150] ^ m[153] ^ m[155] ^ m[157] ^ m[158] ^ m[160] ^ m[162] ^ m[165] ^ m[167] ^ m[169] ^ m[171] ^ m[172] ^ m[175] ^ m[177] ^ m[179] ^ m[180] ^ m[183] ^ m[185] ^ m[187] ^ m[188] ^ m[190] ^ m[192] ^ m[195] ^ m[197] ^ m[199] ^ m[200] ^ m[203] ^ m[205] ^ m[207] ^ m[208] ^ m[210] ^ m[212] ^ m[215] ^ m[217] ^ m[219] ^ m[220] ^ m[222] ^ m[224] ^ m[227] ^ m[229] ^ m[231] ^ m[232] ^ m[234] ^ m[236] ^ m[239] ^ m[241] ^ m[243] ^ m[244] ^ m[247] ^ m[249] ^ m[251] ^ m[253] ^ m[254] ^ m[257] ^ m[259] ^ m[261] ^ m[262] ^ m[265] ^ m[267] ^ m[269] ^ m[270] ^ m[272] ^ m[274] ^ m[277] ^ m[279] ^ m[281] ^ m[283] ^ m[284] ^ m[287] ^ m[289] ^ m[291] ^ m[292] ^ m[295] ^ m[297] ^ m[299] ^ m[300] ^ m[302] ^ m[304] ^ m[307] ^ m[309] ^ m[311] ^ m[312] ^ m[315] ^ m[317] ^ m[319] ^ m[320] ^ m[322] ^ m[324] ^ m[327] ^ m[329] ^ m[331] ^ m[332] ^ m[334] ^ m[336] ^ m[339] ^ m[341] ^ m[343] ^ m[344] ^ m[346] ^ m[348] ^ m[351] ^ m[353] ^ m[354] ^ m[357] ^ m[359] ^ m[361] ^ m[362] ^ m[365] ^ m[367] ^ m[369] ^ m[370] ^ m[372] ^ m[374] ^ m[377] ^ m[379] ^ m[381] ^ m[382] ^ m[385] ^ m[387] ^ m[389] ^ m[390] ^ m[392] ^ m[394] ^ m[397] ^ m[399] ^ m[401] ^ m[402] ^ m[404] ^ m[406] ^ m[409] ^ m[411] ^ m[413] ^ m[414] ^ m[416] ^ m[418] ^ m[421] ^ m[422] ^ m[425] ^ m[427] ^ m[429] ^ m[430] ^ m[432] ^ m[434] ^ m[437] ^ m[439] ^ m[441] ^ m[442] ^ m[444] ^ m[446] ^ m[449] ^ m[451] ^ m[453] ^ m[454] ^ m[456] ^ m[458] ^ m[461] ^ m[462] ^ m[464] ^ m[466] ^ m[469] ^ m[471] ^ m[473] ^ m[474] ^ m[476] ^ m[478] ^ m[481] ^ m[482] ^ m[484] ^ m[486] ^ m[489] ^ m[490] ^ m[492] ^ m[493] ^ m[494] ^ m[496] ^ m[497] ^ m[498] ^ m[499] ^ m[500] ^ m[501];
    assign parity[4] = m[1] ^ m[3] ^ m[5] ^ m[6] ^ m[9] ^ m[11] ^ m[13] ^ m[15] ^ m[17] ^ m[19] ^ m[20] ^ m[23] ^ m[25] ^ m[27] ^ m[29] ^ m[31] ^ m[32] ^ m[35] ^ m[37] ^ m[39] ^ m[41] ^ m[42] ^ m[45] ^ m[47] ^ m[49] ^ m[51] ^ m[52] ^ m[54] ^ m[56] ^ m[58] ^ m[61] ^ m[63] ^ m[65] ^ m[67] ^ m[69] ^ m[71] ^ m[73] ^ m[75] ^ m[76] ^ m[79] ^ m[81] ^ m[83] ^ m[85] ^ m[87] ^ m[88] ^ m[91] ^ m[93] ^ m[95] ^ m[97] ^ m[98] ^ m[101] ^ m[103] ^ m[105] ^ m[107] ^ m[108] ^ m[110] ^ m[112] ^ m[114] ^ m[117] ^ m[119] ^ m[121] ^ m[123] ^ m[125] ^ m[127] ^ m[129] ^ m[130] ^ m[133] ^ m[135] ^ m[137] ^ m[139] ^ m[140] ^ m[143] ^ m[145] ^ m[147] ^ m[149] ^ m[150] ^ m[152] ^ m[154] ^ m[156] ^ m[159] ^ m[161] ^ m[163] ^ m[165] ^ m[167] ^ m[169] ^ m[170] ^ m[173] ^ m[175] ^ m[177] ^ m[179] ^ m[180] ^ m[182] ^ m[184] ^ m[186] ^ m[189] ^ m[191] ^ m[193] ^ m[195] ^ m[197] ^ m[199] ^ m[200] ^ m[202] ^ m[204] ^ m[206] ^ m[209] ^ m[211] ^ m[213] ^ m[215] ^ m[217] ^ m[219] ^ m[220] ^ m[222] ^ m[224] ^ m[226] ^ m[228] ^ m[230] ^ m[233] ^ m[235] ^ m[237] ^ m[239] ^ m[241] ^ m[242] ^ m[245] ^ m[247] ^ m[249] ^ m[251] ^ m[252] ^ m[255] ^ m[257] ^ m[259] ^ m[261] ^ m[262] ^ m[264] ^ m[266] ^ m[268] ^ m[271] ^ m[273] ^ m[275] ^ m[277] ^ m[279] ^ m[281] ^ m[282] ^ m[285] ^ m[287] ^ m[289] ^ m[291] ^ m[292] ^ m[294] ^ m[296] ^ m[298] ^ m[301] ^ m[303] ^ m[305] ^ m[307] ^ m[309] ^ m[311] ^ m[312] ^ m[314] ^ m[316] ^ m[318] ^ m[321] ^ m[323] ^ m[325] ^ m[327] ^ m[329] ^ m[331] ^ m[332] ^ m[334] ^ m[336] ^ m[338] ^ m[340] ^ m[342] ^ m[345] ^ m[347] ^ m[349] ^ m[351] ^ m[352] ^ m[355] ^ m[357] ^ m[359] ^ m[361] ^ m[362] ^ m[364] ^ m[366] ^ m[368] ^ m[371] ^ m[373] ^ m[375] ^ m[377] ^ m[379] ^ m[381] ^ m[382] ^ m[384] ^ m[386] ^ m[388] ^ m[391] ^ m[393] ^ m[395] ^ m[397] ^ m[399] ^ m[401] ^ m[402] ^ m[404] ^ m[406] ^ m[408] ^ m[410] ^ m[412] ^ m[415] ^ m[417] ^ m[419] ^ m[421] ^ m[422] ^ m[424] ^ m[426] ^ m[428] ^ m[431] ^ m[433] ^ m[435] ^ m[437] ^ m[439] ^ m[441] ^ m[442] ^ m[444] ^ m[446] ^ m[448] ^ m[450] ^ m[452] ^ m[455] ^ m[457] ^ m[459] ^ m[461] ^ m[462] ^ m[464] ^ m[466] ^ m[468] ^ m[470] ^ m[472] ^ m[475] ^ m[477] ^ m[479] ^ m[481] ^ m[482] ^ m[484] ^ m[486] ^ m[488] ^ m[491] ^ m[492] ^ m[493] ^ m[494] ^ m[495] ^ m[497] ^ m[498] ^ m[499] ^ m[500] ^ m[501];
    assign parity[5] = m[1] ^ m[3] ^ m[4] ^ m[7] ^ m[9] ^ m[11] ^ m[13] ^ m[15] ^ m[17] ^ m[18] ^ m[21] ^ m[23] ^ m[25] ^ m[27] ^ m[29] ^ m[30] ^ m[33] ^ m[35] ^ m[37] ^ m[39] ^ m[41] ^ m[42] ^ m[44] ^ m[46] ^ m[48] ^ m[50] ^ m[53] ^ m[55] ^ m[57] ^ m[59] ^ m[61] ^ m[63] ^ m[65] ^ m[67] ^ m[69] ^ m[71] ^ m[73] ^ m[74] ^ m[77] ^ m[79] ^ m[81] ^ m[83] ^ m[85] ^ m[86] ^ m[89] ^ m[91] ^ m[93] ^ m[95] ^ m[97] ^ m[98] ^ m[100] ^ m[102] ^ m[104] ^ m[106] ^ m[109] ^ m[111] ^ m[113] ^ m[115] ^ m[117] ^ m[119] ^ m[121] ^ m[123] ^ m[125] ^ m[127] ^ m[128] ^ m[131] ^ m[133] ^ m[135] ^ m[137] ^ m[139] ^ m[140] ^ m[142] ^ m[144] ^ m[146] ^ m[148] ^ m[151] ^ m[153] ^ m[155] ^ m[157] ^ m[159] ^ m[161] ^ m[163] ^ m[165] ^ m[167] ^ m[169] ^ m[170] ^ m[172] ^ m[174] ^ m[176] ^ m[178] ^ m[181] ^ m[183] ^ m[185] ^ m[187] ^ m[189] ^ m[191] ^ m[193] ^ m[195] ^ m[197] ^ m[199] ^ m[200] ^ m[202] ^ m[204] ^ m[206] ^ m[208] ^ m[210] ^ m[212] ^ m[214] ^ m[216] ^ m[218] ^ m[221] ^ m[223] ^ m[225] ^ m[227] ^ m[229] ^ m[231] ^ m[233] ^ m[235] ^ m[237] ^ m[239] ^ m[240] ^ m[243] ^ m[245] ^ m[247] ^ m[249] ^ m[251] ^ m[252] ^ m[254] ^ m[256] ^ m[258] ^ m[260] ^ m[263] ^ m[265] ^ m[267] ^ m[269] ^ m[271] ^ m[273] ^ m[275] ^ m[277] ^ m[279] ^ m[281] ^ m[282] ^ m[284] ^ m[286] ^ m[288] ^ m[290] ^ m[293] ^ m[295] ^ m[297] ^ m[299] ^ m[301] ^ m[303] ^ m[305] ^ m[307] ^ m[309] ^ m[311] ^ m[312] ^ m[314] ^ m[316] ^ m[318] ^ m[320] ^ m[322] ^ m[324] ^ m[326] ^ m[328] ^ m[330] ^ m[333] ^ m[335] ^ m[337] ^ m[339] ^ m[341] ^ m[343] ^ m[345] ^ m[347] ^ m[349] ^ m[351] ^ m[352] ^ m[354] ^ m[356] ^ m[358] ^ m[360] ^ m[363] ^ m[365] ^ m[367] ^ m[369] ^ m[371] ^ m[373] ^ m[375] ^ m[377] ^ m[379] ^ m[381] ^ m[382] ^ m[384] ^ m[386] ^ m[388] ^ m[390] ^ m[392] ^ m[394] ^ m[396] ^ m[398] ^ m[400] ^ m[403] ^ m[405] ^ m[407] ^ m[409] ^ m[411] ^ m[413] ^ m[415] ^ m[417] ^ m[419] ^ m[421] ^ m[422] ^ m[424] ^ m[426] ^ m[428] ^ m[430] ^ m[432] ^ m[434] ^ m[436] ^ m[438] ^ m[440] ^ m[443] ^ m[445] ^ m[447] ^ m[449] ^ m[451] ^ m[453] ^ m[455] ^ m[457] ^ m[459] ^ m[461] ^ m[462] ^ m[464] ^ m[466] ^ m[468] ^ m[470] ^ m[472] ^ m[474] ^ m[476] ^ m[478] ^ m[480] ^ m[483] ^ m[485] ^ m[487] ^ m[489] ^ m[491] ^ m[492] ^ m[493] ^ m[494] ^ m[495] ^ m[496] ^ m[498] ^ m[499] ^ m[500] ^ m[501];
    assign parity[6] = m[1] ^ m[2] ^ m[5] ^ m[7] ^ m[9] ^ m[11] ^ m[13] ^ m[15] ^ m[16] ^ m[19] ^ m[21] ^ m[23] ^ m[25] ^ m[27] ^ m[29] ^ m[30] ^ m[32] ^ m[34] ^ m[36] ^ m[38] ^ m[40] ^ m[43] ^ m[45] ^ m[47] ^ m[49] ^ m[51] ^ m[53] ^ m[55] ^ m[57] ^ m[59] ^ m[61] ^ m[63] ^ m[65] ^ m[67] ^ m[69] ^ m[71] ^ m[72] ^ m[75] ^ m[77] ^ m[79] ^ m[81] ^ m[83] ^ m[85] ^ m[86] ^ m[88] ^ m[90] ^ m[92] ^ m[94] ^ m[96] ^ m[99] ^ m[101] ^ m[103] ^ m[105] ^ m[107] ^ m[109] ^ m[111] ^ m[113] ^ m[115] ^ m[117] ^ m[119] ^ m[121] ^ m[123] ^ m[125] ^ m[127] ^ m[128] ^ m[130] ^ m[132] ^ m[134] ^ m[136] ^ m[138] ^ m[141] ^ m[143] ^ m[145] ^ m[147] ^ m[149] ^ m[151] ^ m[153] ^ m[155] ^ m[157] ^ m[159] ^ m[161] ^ m[163] ^ m[165] ^ m[167] ^ m[169] ^ m[170] ^ m[172] ^ m[174] ^ m[176] ^ m[178] ^ m[180] ^ m[182] ^ m[184] ^ m[186] ^ m[188] ^ m[190] ^ m[192] ^ m[194] ^ m[196] ^ m[198] ^ m[201] ^ m[203] ^ m[205] ^ m[207] ^ m[209] ^ m[211] ^ m[213] ^ m[215] ^ m[217] ^ m[219] ^ m[221] ^ m[223] ^ m[225] ^ m[227] ^ m[229] ^ m[231] ^ m[233] ^ m[235] ^ m[237] ^ m[239] ^ m[240] ^ m[242] ^ m[244] ^ m[246] ^ m[248] ^ m[250] ^ m[253] ^ m[255] ^ m[257] ^ m[259] ^ m[261] ^ m[263] ^ m[265] ^ m[267] ^ m[269] ^ m[271] ^ m[273] ^ m[275] ^ m[277] ^ m[279] ^ m[281] ^ m[282] ^ m[284] ^ m[286] ^ m[288] ^ m[290] ^ m[292] ^ m[294] ^ m[296] ^ m[298] ^ m[300] ^ m[302] ^ m[304] ^ m[306] ^ m[308] ^ m[310] ^ m[313] ^ m[315] ^ m[317] ^ m[319] ^ m[321] ^ m[323] ^ m[325] ^ m[327] ^ m[329] ^ m[331] ^ m[333] ^ m[335] ^ m[337] ^ m[339] ^ m[341] ^ m[343] ^ m[345] ^ m[347] ^ m[349] ^ m[351] ^ m[352] ^ m[354] ^ m[356] ^ m[358] ^ m[360] ^ m[362] ^ m[364] ^ m[366] ^ m[368] ^ m[370] ^ m[372] ^ m[374] ^ m[376] ^ m[378] ^ m[380] ^ m[383] ^ m[385] ^ m[387] ^ m[389] ^ m[391] ^ m[393] ^ m[395] ^ m[397] ^ m[399] ^ m[401] ^ m[403] ^ m[405] ^ m[407] ^ m[409] ^ m[411] ^ m[413] ^ m[415] ^ m[417] ^ m[419] ^ m[421] ^ m[422] ^ m[424] ^ m[426] ^ m[428] ^ m[430] ^ m[432] ^ m[434] ^ m[436] ^ m[438] ^ m[440] ^ m[442] ^ m[444] ^ m[446] ^ m[448] ^ m[450] ^ m[452] ^ m[454] ^ m[456] ^ m[458] ^ m[460] ^ m[463] ^ m[465] ^ m[467] ^ m[469] ^ m[471] ^ m[473] ^ m[475] ^ m[477] ^ m[479] ^ m[481] ^ m[483] ^ m[485] ^ m[487] ^ m[489] ^ m[491] ^ m[492] ^ m[493] ^ m[494] ^ m[495] ^ m[496] ^ m[497] ^ m[499] ^ m[500] ^ m[501];
    assign parity[7] = m[0] ^ m[3] ^ m[5] ^ m[7] ^ m[9] ^ m[11] ^ m[13] ^ m[15] ^ m[16] ^ m[18] ^ m[20] ^ m[22] ^ m[24] ^ m[26] ^ m[28] ^ m[31] ^ m[33] ^ m[35] ^ m[37] ^ m[39] ^ m[41] ^ m[43] ^ m[45] ^ m[47] ^ m[49] ^ m[51] ^ m[53] ^ m[55] ^ m[57] ^ m[59] ^ m[61] ^ m[63] ^ m[65] ^ m[67] ^ m[69] ^ m[71] ^ m[72] ^ m[74] ^ m[76] ^ m[78] ^ m[80] ^ m[82] ^ m[84] ^ m[87] ^ m[89] ^ m[91] ^ m[93] ^ m[95] ^ m[97] ^ m[99] ^ m[101] ^ m[103] ^ m[105] ^ m[107] ^ m[109] ^ m[111] ^ m[113] ^ m[115] ^ m[117] ^ m[119] ^ m[121] ^ m[123] ^ m[125] ^ m[127] ^ m[128] ^ m[130] ^ m[132] ^ m[134] ^ m[136] ^ m[138] ^ m[140] ^ m[142] ^ m[144] ^ m[146] ^ m[148] ^ m[150] ^ m[152] ^ m[154] ^ m[156] ^ m[158] ^ m[160] ^ m[162] ^ m[164] ^ m[166] ^ m[168] ^ m[171] ^ m[173] ^ m[175] ^ m[177] ^ m[179] ^ m[181] ^ m[183] ^ m[185] ^ m[187] ^ m[189] ^ m[191] ^ m[193] ^ m[195] ^ m[197] ^ m[199] ^ m[201] ^ m[203] ^ m[205] ^ m[207] ^ m[209] ^ m[211] ^ m[213] ^ m[215] ^ m[217] ^ m[219] ^ m[221] ^ m[223] ^ m[225] ^ m[227] ^ m[229] ^ m[231] ^ m[233] ^ m[235] ^ m[237] ^ m[239] ^ m[240] ^ m[242] ^ m[244] ^ m[246] ^ m[248] ^ m[250] ^ m[252] ^ m[254] ^ m[256] ^ m[258] ^ m[260] ^ m[262] ^ m[264] ^ m[266] ^ m[268] ^ m[270] ^ m[272] ^ m[274] ^ m[276] ^ m[278] ^ m[280] ^ m[283] ^ m[285] ^ m[287] ^ m[289] ^ m[291] ^ m[293] ^ m[295] ^ m[297] ^ m[299] ^ m[301] ^ m[303] ^ m[305] ^ m[307] ^ m[309] ^ m[311] ^ m[313] ^ m[315] ^ m[317] ^ m[319] ^ m[321] ^ m[323] ^ m[325] ^ m[327] ^ m[329] ^ m[331] ^ m[333] ^ m[335] ^ m[337] ^ m[339] ^ m[341] ^ m[343] ^ m[345] ^ m[347] ^ m[349] ^ m[351] ^ m[352] ^ m[354] ^ m[356] ^ m[358] ^ m[360] ^ m[362] ^ m[364] ^ m[366] ^ m[368] ^ m[370] ^ m[372] ^ m[374] ^ m[376] ^ m[378] ^ m[380] ^ m[382] ^ m[384] ^ m[386] ^ m[388] ^ m[390] ^ m[392] ^ m[394] ^ m[396] ^ m[398] ^ m[400] ^ m[402] ^ m[404] ^ m[406] ^ m[408] ^ m[410] ^ m[412] ^ m[414] ^ m[416] ^ m[418] ^ m[420] ^ m[423] ^ m[425] ^ m[427] ^ m[429] ^ m[431] ^ m[433] ^ m[435] ^ m[437] ^ m[439] ^ m[441] ^ m[443] ^ m[445] ^ m[447] ^ m[449] ^ m[451] ^ m[453] ^ m[455] ^ m[457] ^ m[459] ^ m[461] ^ m[463] ^ m[465] ^ m[467] ^ m[469] ^ m[471] ^ m[473] ^ m[475] ^ m[477] ^ m[479] ^ m[481] ^ m[483] ^ m[485] ^ m[487] ^ m[489] ^ m[491] ^ m[492] ^ m[493] ^ m[494] ^ m[495] ^ m[496] ^ m[497] ^ m[498] ^ m[500] ^ m[501];
    assign parity[8] = m[0] ^ m[2] ^ m[4] ^ m[6] ^ m[8] ^ m[10] ^ m[12] ^ m[14] ^ m[17] ^ m[19] ^ m[21] ^ m[23] ^ m[25] ^ m[27] ^ m[29] ^ m[31] ^ m[33] ^ m[35] ^ m[37] ^ m[39] ^ m[41] ^ m[43] ^ m[45] ^ m[47] ^ m[49] ^ m[51] ^ m[53] ^ m[55] ^ m[57] ^ m[59] ^ m[61] ^ m[63] ^ m[65] ^ m[67] ^ m[69] ^ m[71] ^ m[72] ^ m[74] ^ m[76] ^ m[78] ^ m[80] ^ m[82] ^ m[84] ^ m[86] ^ m[88] ^ m[90] ^ m[92] ^ m[94] ^ m[96] ^ m[98] ^ m[100] ^ m[102] ^ m[104] ^ m[106] ^ m[108] ^ m[110] ^ m[112] ^ m[114] ^ m[116] ^ m[118] ^ m[120] ^ m[122] ^ m[124] ^ m[126] ^ m[129] ^ m[131] ^ m[133] ^ m[135] ^ m[137] ^ m[139] ^ m[141] ^ m[143] ^ m[145] ^ m[147] ^ m[149] ^ m[151] ^ m[153] ^ m[155] ^ m[157] ^ m[159] ^ m[161] ^ m[163] ^ m[165] ^ m[167] ^ m[169] ^ m[171] ^ m[173] ^ m[175] ^ m[177] ^ m[179] ^ m[181] ^ m[183] ^ m[185] ^ m[187] ^ m[189] ^ m[191] ^ m[193] ^ m[195] ^ m[197] ^ m[199] ^ m[201] ^ m[203] ^ m[205] ^ m[207] ^ m[209] ^ m[211] ^ m[213] ^ m[215] ^ m[217] ^ m[219] ^ m[221] ^ m[223] ^ m[225] ^ m[227] ^ m[229] ^ m[231] ^ m[233] ^ m[235] ^ m[237] ^ m[239] ^ m[240] ^ m[242] ^ m[244] ^ m[246] ^ m[248] ^ m[250] ^ m[252] ^ m[254] ^ m[256] ^ m[258] ^ m[260] ^ m[262] ^ m[264] ^ m[266] ^ m[268] ^ m[270] ^ m[272] ^ m[274] ^ m[276] ^ m[278] ^ m[280] ^ m[282] ^ m[284] ^ m[286] ^ m[288] ^ m[290] ^ m[292] ^ m[294] ^ m[296] ^ m[298] ^ m[300] ^ m[302] ^ m[304] ^ m[306] ^ m[308] ^ m[310] ^ m[312] ^ m[314] ^ m[316] ^ m[318] ^ m[320] ^ m[322] ^ m[324] ^ m[326] ^ m[328] ^ m[330] ^ m[332] ^ m[334] ^ m[336] ^ m[338] ^ m[340] ^ m[342] ^ m[344] ^ m[346] ^ m[348] ^ m[350] ^ m[353] ^ m[355] ^ m[357] ^ m[359] ^ m[361] ^ m[363] ^ m[365] ^ m[367] ^ m[369] ^ m[371] ^ m[373] ^ m[375] ^ m[377] ^ m[379] ^ m[381] ^ m[383] ^ m[385] ^ m[387] ^ m[389] ^ m[391] ^ m[393] ^ m[395] ^ m[397] ^ m[399] ^ m[401] ^ m[403] ^ m[405] ^ m[407] ^ m[409] ^ m[411] ^ m[413] ^ m[415] ^ m[417] ^ m[419] ^ m[421] ^ m[423] ^ m[425] ^ m[427] ^ m[429] ^ m[431] ^ m[433] ^ m[435] ^ m[437] ^ m[439] ^ m[441] ^ m[443] ^ m[445] ^ m[447] ^ m[449] ^ m[451] ^ m[453] ^ m[455] ^ m[457] ^ m[459] ^ m[461] ^ m[463] ^ m[465] ^ m[467] ^ m[469] ^ m[471] ^ m[473] ^ m[475] ^ m[477] ^ m[479] ^ m[481] ^ m[483] ^ m[485] ^ m[487] ^ m[489] ^ m[491] ^ m[492] ^ m[493] ^ m[494] ^ m[495] ^ m[496] ^ m[497] ^ m[498] ^ m[499] ^ m[501];
    assign parity[9] = m[0] ^ m[2] ^ m[4] ^ m[6] ^ m[8] ^ m[10] ^ m[12] ^ m[14] ^ m[16] ^ m[18] ^ m[20] ^ m[22] ^ m[24] ^ m[26] ^ m[28] ^ m[30] ^ m[32] ^ m[34] ^ m[36] ^ m[38] ^ m[40] ^ m[42] ^ m[44] ^ m[46] ^ m[48] ^ m[50] ^ m[52] ^ m[54] ^ m[56] ^ m[58] ^ m[60] ^ m[62] ^ m[64] ^ m[66] ^ m[68] ^ m[70] ^ m[73] ^ m[75] ^ m[77] ^ m[79] ^ m[81] ^ m[83] ^ m[85] ^ m[87] ^ m[89] ^ m[91] ^ m[93] ^ m[95] ^ m[97] ^ m[99] ^ m[101] ^ m[103] ^ m[105] ^ m[107] ^ m[109] ^ m[111] ^ m[113] ^ m[115] ^ m[117] ^ m[119] ^ m[121] ^ m[123] ^ m[125] ^ m[127] ^ m[129] ^ m[131] ^ m[133] ^ m[135] ^ m[137] ^ m[139] ^ m[141] ^ m[143] ^ m[145] ^ m[147] ^ m[149] ^ m[151] ^ m[153] ^ m[155] ^ m[157] ^ m[159] ^ m[161] ^ m[163] ^ m[165] ^ m[167] ^ m[169] ^ m[171] ^ m[173] ^ m[175] ^ m[177] ^ m[179] ^ m[181] ^ m[183] ^ m[185] ^ m[187] ^ m[189] ^ m[191] ^ m[193] ^ m[195] ^ m[197] ^ m[199] ^ m[201] ^ m[203] ^ m[205] ^ m[207] ^ m[209] ^ m[211] ^ m[213] ^ m[215] ^ m[217] ^ m[219] ^ m[221] ^ m[223] ^ m[225] ^ m[227] ^ m[229] ^ m[231] ^ m[233] ^ m[235] ^ m[237] ^ m[239] ^ m[240] ^ m[242] ^ m[244] ^ m[246] ^ m[248] ^ m[250] ^ m[252] ^ m[254] ^ m[256] ^ m[258] ^ m[260] ^ m[262] ^ m[264] ^ m[266] ^ m[268] ^ m[270] ^ m[272] ^ m[274] ^ m[276] ^ m[278] ^ m[280] ^ m[282] ^ m[284] ^ m[286] ^ m[288] ^ m[290] ^ m[292] ^ m[294] ^ m[296] ^ m[298] ^ m[300] ^ m[302] ^ m[304] ^ m[306] ^ m[308] ^ m[310] ^ m[312] ^ m[314] ^ m[316] ^ m[318] ^ m[320] ^ m[322] ^ m[324] ^ m[326] ^ m[328] ^ m[330] ^ m[332] ^ m[334] ^ m[336] ^ m[338] ^ m[340] ^ m[342] ^ m[344] ^ m[346] ^ m[348] ^ m[350] ^ m[352] ^ m[354] ^ m[356] ^ m[358] ^ m[360] ^ m[362] ^ m[364] ^ m[366] ^ m[368] ^ m[370] ^ m[372] ^ m[374] ^ m[376] ^ m[378] ^ m[380] ^ m[382] ^ m[384] ^ m[386] ^ m[388] ^ m[390] ^ m[392] ^ m[394] ^ m[396] ^ m[398] ^ m[400] ^ m[402] ^ m[404] ^ m[406] ^ m[408] ^ m[410] ^ m[412] ^ m[414] ^ m[416] ^ m[418] ^ m[420] ^ m[422] ^ m[424] ^ m[426] ^ m[428] ^ m[430] ^ m[432] ^ m[434] ^ m[436] ^ m[438] ^ m[440] ^ m[442] ^ m[444] ^ m[446] ^ m[448] ^ m[450] ^ m[452] ^ m[454] ^ m[456] ^ m[458] ^ m[460] ^ m[462] ^ m[464] ^ m[466] ^ m[468] ^ m[470] ^ m[472] ^ m[474] ^ m[476] ^ m[478] ^ m[480] ^ m[482] ^ m[484] ^ m[486] ^ m[488] ^ m[490] ^ m[492] ^ m[493] ^ m[494] ^ m[495] ^ m[496] ^ m[497] ^ m[498] ^ m[499] ^ m[500];
  end else if ((CodewordWidth == 1024) && (MessageWidth == 1013)) begin : gen_1024_1013
    `BR_ASSERT_STATIC(parity_width_matches_a, ParityWidth == 11)
    assign parity[0] = m[0] ^ m[2] ^ m[4] ^ m[6] ^ m[8] ^ m[10] ^ m[12] ^ m[14] ^ m[16] ^ m[18] ^ m[20] ^ m[22] ^ m[24] ^ m[26] ^ m[28] ^ m[30] ^ m[31] ^ m[33] ^ m[36] ^ m[38] ^ m[40] ^ m[42] ^ m[44] ^ m[46] ^ m[48] ^ m[50] ^ m[52] ^ m[54] ^ m[56] ^ m[58] ^ m[59] ^ m[62] ^ m[64] ^ m[65] ^ m[68] ^ m[70] ^ m[72] ^ m[74] ^ m[76] ^ m[78] ^ m[80] ^ m[82] ^ m[83] ^ m[86] ^ m[88] ^ m[90] ^ m[92] ^ m[93] ^ m[96] ^ m[98] ^ m[100] ^ m[102] ^ m[103] ^ m[106] ^ m[108] ^ m[110] ^ m[112] ^ m[114] ^ m[116] ^ m[117] ^ m[119] ^ m[122] ^ m[124] ^ m[126] ^ m[128] ^ m[130] ^ m[131] ^ m[134] ^ m[136] ^ m[137] ^ m[139] ^ m[142] ^ m[143] ^ m[146] ^ m[148] ^ m[150] ^ m[152] ^ m[153] ^ m[156] ^ m[158] ^ m[160] ^ m[162] ^ m[164] ^ m[165] ^ m[168] ^ m[170] ^ m[171] ^ m[173] ^ m[176] ^ m[177] ^ m[180] ^ m[183] ^ m[186] ^ m[189] ^ m[190] ^ m[195] ^ m[197] ^ m[199] ^ m[202] ^ m[203] ^ m[206] ^ m[209] ^ m[211] ^ m[212] ^ m[216] ^ m[217] ^ m[222] ^ m[225] ^ m[227] ^ m[229] ^ m[232] ^ m[233] ^ m[235] ^ m[237] ^ m[241] ^ m[244] ^ m[246] ^ m[248] ^ m[252] ^ m[253] ^ m[256] ^ m[260] ^ m[262] ^ m[263] ^ m[268] ^ m[270] ^ m[272] ^ m[276] ^ m[278] ^ m[281] ^ m[282] ^ m[285] ^ m[288] ^ m[290] ^ m[294] ^ m[295] ^ m[296] ^ m[299] ^ m[302] ^ m[303] ^ m[306] ^ m[308] ^ m[311] ^ m[313] ^ m[315] ^ m[317] ^ m[319] ^ m[321] ^ m[323] ^ m[325] ^ m[326] ^ m[329] ^ m[331] ^ m[332] ^ m[335] ^ m[337] ^ m[339] ^ m[341] ^ m[343] ^ m[345] ^ m[346] ^ m[349] ^ m[351] ^ m[352] ^ m[355] ^ m[357] ^ m[359] ^ m[361] ^ m[362] ^ m[365] ^ m[367] ^ m[368] ^ m[371] ^ m[373] ^ m[374] ^ m[377] ^ m[379] ^ m[380] ^ m[382] ^ m[385] ^ m[386] ^ m[388] ^ m[391] ^ m[392] ^ m[395] ^ m[397] ^ m[399] ^ m[401] ^ m[403] ^ m[405] ^ m[407] ^ m[409] ^ m[410] ^ m[412] ^ m[415] ^ m[417] ^ m[419] ^ m[421] ^ m[423] ^ m[425] ^ m[427] ^ m[428] ^ m[431] ^ m[433] ^ m[434] ^ m[437] ^ m[439] ^ m[440] ^ m[442] ^ m[445] ^ m[447] ^ m[448] ^ m[450] ^ m[452] ^ m[454] ^ m[457] ^ m[459] ^ m[461] ^ m[463] ^ m[465] ^ m[467] ^ m[468] ^ m[471] ^ m[473] ^ m[475] ^ m[477] ^ m[478] ^ m[480] ^ m[483] ^ m[485] ^ m[486] ^ m[488] ^ m[491] ^ m[492] ^ m[494] ^ m[497] ^ m[499] ^ m[501] ^ m[503] ^ m[504] ^ m[507] ^ m[509] ^ m[510] ^ m[512] ^ m[515] ^ m[516] ^ m[519] ^ m[521] ^ m[523] ^ m[524] ^ m[526] ^ m[528] ^ m[530] ^ m[532] ^ m[535] ^ m[537] ^ m[539] ^ m[541] ^ m[542] ^ m[545] ^ m[547] ^ m[549] ^ m[550] ^ m[552] ^ m[554] ^ m[557] ^ m[558] ^ m[560] ^ m[562] ^ m[564] ^ m[566] ^ m[568] ^ m[570] ^ m[572] ^ m[574] ^ m[575] ^ m[578] ^ m[580] ^ m[581] ^ m[584] ^ m[586] ^ m[588] ^ m[590] ^ m[592] ^ m[593] ^ m[595] ^ m[598] ^ m[600] ^ m[601] ^ m[604] ^ m[605] ^ m[608] ^ m[610] ^ m[611] ^ m[614] ^ m[616] ^ m[618] ^ m[620] ^ m[622] ^ m[623] ^ m[625] ^ m[628] ^ m[630] ^ m[631] ^ m[633] ^ m[635] ^ m[638] ^ m[640] ^ m[642] ^ m[644] ^ m[645] ^ m[648] ^ m[650] ^ m[652] ^ m[653] ^ m[655] ^ m[658] ^ m[660] ^ m[661] ^ m[664] ^ m[666] ^ m[668] ^ m[670] ^ m[671] ^ m[673] ^ m[676] ^ m[678] ^ m[680] ^ m[681] ^ m[683] ^ m[685] ^ m[688] ^ m[690] ^ m[691] ^ m[693] ^ m[695] ^ m[697] ^ m[700] ^ m[702] ^ m[704] ^ m[705] ^ m[708] ^ m[710] ^ m[711] ^ m[714] ^ m[716] ^ m[718] ^ m[720] ^ m[721] ^ m[723] ^ m[726] ^ m[728] ^ m[730] ^ m[731] ^ m[733] ^ m[735] ^ m[738] ^ m[740] ^ m[741] ^ m[744] ^ m[745] ^ m[747] ^ m[750] ^ m[752] ^ m[754] ^ m[755] ^ m[757] ^ m[759] ^ m[762] ^ m[764] ^ m[765] ^ m[767] ^ m[769] ^ m[771] ^ m[774] ^ m[775] ^ m[777] ^ m[780] ^ m[781] ^ m[783] ^ m[785] ^ m[788] ^ m[790] ^ m[792] ^ m[794] ^ m[795] ^ m[797] ^ m[800] ^ m[802] ^ m[803] ^ m[805] ^ m[807] ^ m[809] ^ m[812] ^ m[814] ^ m[816] ^ m[818] ^ m[819] ^ m[821] ^ m[822] ^ m[825] ^ m[827] ^ m[829] ^ m[830] ^ m[832] ^ m[834] ^ m[836] ^ m[837] ^ m[839] ^ m[841] ^ m[843] ^ m[845] ^ m[846] ^ m[847] ^ m[849] ^ m[852] ^ m[853] ^ m[855] ^ m[856] ^ m[859] ^ m[860] ^ m[862] ^ m[864] ^ m[865] ^ m[866] ^ m[869] ^ m[870] ^ m[872] ^ m[875] ^ m[877] ^ m[878] ^ m[880] ^ m[881] ^ m[882] ^ m[884] ^ m[886] ^ m[887] ^ m[889] ^ m[892] ^ m[893] ^ m[895] ^ m[896] ^ m[898] ^ m[899] ^ m[901] ^ m[902] ^ m[906] ^ m[907] ^ m[908] ^ m[911] ^ m[912] ^ m[915] ^ m[916] ^ m[917] ^ m[919] ^ m[922] ^ m[924] ^ m[926] ^ m[927] ^ m[928] ^ m[931] ^ m[933] ^ m[934] ^ m[936] ^ m[938] ^ m[940] ^ m[942] ^ m[943] ^ m[945] ^ m[947] ^ m[948] ^ m[950] ^ m[951] ^ m[953] ^ m[955] ^ m[957] ^ m[958] ^ m[960] ^ m[963] ^ m[964] ^ m[966] ^ m[967] ^ m[968] ^ m[970] ^ m[972] ^ m[973] ^ m[975] ^ m[976] ^ m[978] ^ m[979] ^ m[982] ^ m[983] ^ m[984] ^ m[986] ^ m[988] ^ m[990] ^ m[991] ^ m[993] ^ m[995] ^ m[996] ^ m[997] ^ m[1000] ^ m[1001] ^ m[1002] ^ m[1004] ^ m[1005] ^ m[1006] ^ m[1008] ^ m[1009] ^ m[1011] ^ m[1012];
    assign parity[1] = m[0] ^ m[2] ^ m[4] ^ m[6] ^ m[8] ^ m[10] ^ m[12] ^ m[14] ^ m[16] ^ m[18] ^ m[20] ^ m[22] ^ m[24] ^ m[26] ^ m[27] ^ m[29] ^ m[32] ^ m[34] ^ m[36] ^ m[38] ^ m[40] ^ m[42] ^ m[44] ^ m[46] ^ m[48] ^ m[50] ^ m[52] ^ m[54] ^ m[55] ^ m[58] ^ m[60] ^ m[61] ^ m[64] ^ m[66] ^ m[68] ^ m[70] ^ m[72] ^ m[74] ^ m[76] ^ m[78] ^ m[79] ^ m[82] ^ m[84] ^ m[86] ^ m[88] ^ m[89] ^ m[92] ^ m[94] ^ m[96] ^ m[98] ^ m[99] ^ m[102] ^ m[104] ^ m[106] ^ m[108] ^ m[110] ^ m[112] ^ m[113] ^ m[115] ^ m[118] ^ m[120] ^ m[122] ^ m[124] ^ m[126] ^ m[127] ^ m[130] ^ m[132] ^ m[133] ^ m[135] ^ m[138] ^ m[140] ^ m[142] ^ m[143] ^ m[146] ^ m[148] ^ m[149] ^ m[152] ^ m[154] ^ m[156] ^ m[158] ^ m[160] ^ m[161] ^ m[164] ^ m[166] ^ m[167] ^ m[169] ^ m[172] ^ m[174] ^ m[176] ^ m[177] ^ m[180] ^ m[183] ^ m[186] ^ m[187] ^ m[191] ^ m[195] ^ m[197] ^ m[199] ^ m[202] ^ m[204] ^ m[206] ^ m[208] ^ m[211] ^ m[213] ^ m[214] ^ m[219] ^ m[221] ^ m[224] ^ m[227] ^ m[228] ^ m[230] ^ m[234] ^ m[236] ^ m[238] ^ m[241] ^ m[243] ^ m[247] ^ m[249] ^ m[250] ^ m[254] ^ m[256] ^ m[260] ^ m[262] ^ m[265] ^ m[267] ^ m[269] ^ m[273] ^ m[275] ^ m[279] ^ m[280] ^ m[283] ^ m[285] ^ m[288] ^ m[291] ^ m[292] ^ m[295] ^ m[298] ^ m[299] ^ m[301] ^ m[305] ^ m[306] ^ m[308] ^ m[311] ^ m[313] ^ m[315] ^ m[317] ^ m[319] ^ m[321] ^ m[322] ^ m[325] ^ m[327] ^ m[328] ^ m[331] ^ m[333] ^ m[335] ^ m[337] ^ m[339] ^ m[341] ^ m[342] ^ m[345] ^ m[347] ^ m[348] ^ m[351] ^ m[353] ^ m[355] ^ m[357] ^ m[358] ^ m[361] ^ m[363] ^ m[364] ^ m[367] ^ m[369] ^ m[370] ^ m[373] ^ m[375] ^ m[376] ^ m[378] ^ m[381] ^ m[383] ^ m[384] ^ m[386] ^ m[389] ^ m[391] ^ m[392] ^ m[395] ^ m[397] ^ m[399] ^ m[401] ^ m[403] ^ m[405] ^ m[406] ^ m[408] ^ m[411] ^ m[413] ^ m[415] ^ m[417] ^ m[419] ^ m[421] ^ m[422] ^ m[424] ^ m[427] ^ m[429] ^ m[431] ^ m[433] ^ m[435] ^ m[436] ^ m[438] ^ m[441] ^ m[443] ^ m[444] ^ m[446] ^ m[449] ^ m[451] ^ m[452] ^ m[454] ^ m[457] ^ m[459] ^ m[461] ^ m[463] ^ m[464] ^ m[467] ^ m[469] ^ m[471] ^ m[473] ^ m[474] ^ m[476] ^ m[479] ^ m[481] ^ m[483] ^ m[484] ^ m[487] ^ m[489] ^ m[490] ^ m[492] ^ m[494] ^ m[497] ^ m[499] ^ m[500] ^ m[503] ^ m[505] ^ m[506] ^ m[508] ^ m[511] ^ m[513] ^ m[515] ^ m[516] ^ m[518] ^ m[520] ^ m[522] ^ m[525] ^ m[527] ^ m[528] ^ m[530] ^ m[532] ^ m[534] ^ m[537] ^ m[538] ^ m[541] ^ m[543] ^ m[545] ^ m[546] ^ m[548] ^ m[551] ^ m[553] ^ m[554] ^ m[557] ^ m[558] ^ m[560] ^ m[562] ^ m[564] ^ m[566] ^ m[568] ^ m[570] ^ m[571] ^ m[573] ^ m[576] ^ m[578] ^ m[580] ^ m[582] ^ m[584] ^ m[586] ^ m[588] ^ m[589] ^ m[591] ^ m[594] ^ m[596] ^ m[597] ^ m[600] ^ m[602] ^ m[604] ^ m[605] ^ m[607] ^ m[610] ^ m[612] ^ m[613] ^ m[616] ^ m[618] ^ m[619] ^ m[622] ^ m[624] ^ m[626] ^ m[627] ^ m[629] ^ m[632] ^ m[634] ^ m[635] ^ m[638] ^ m[640] ^ m[641] ^ m[644] ^ m[646] ^ m[648] ^ m[649] ^ m[651] ^ m[654] ^ m[656] ^ m[658] ^ m[660] ^ m[661] ^ m[664] ^ m[666] ^ m[667] ^ m[669] ^ m[672] ^ m[674] ^ m[676] ^ m[677] ^ m[679] ^ m[682] ^ m[684] ^ m[685] ^ m[687] ^ m[689] ^ m[692] ^ m[694] ^ m[695] ^ m[697] ^ m[700] ^ m[702] ^ m[704] ^ m[705] ^ m[707] ^ m[710] ^ m[712] ^ m[714] ^ m[716] ^ m[717] ^ m[719] ^ m[722] ^ m[724] ^ m[726] ^ m[727] ^ m[729] ^ m[732] ^ m[734] ^ m[735] ^ m[737] ^ m[740] ^ m[742] ^ m[743] ^ m[745] ^ m[748] ^ m[750] ^ m[751] ^ m[753] ^ m[756] ^ m[758] ^ m[759] ^ m[761] ^ m[763] ^ m[766] ^ m[768] ^ m[769] ^ m[771] ^ m[773] ^ m[775] ^ m[778] ^ m[779] ^ m[781] ^ m[784] ^ m[785] ^ m[788] ^ m[790] ^ m[791] ^ m[793] ^ m[796] ^ m[798] ^ m[799] ^ m[801] ^ m[804] ^ m[806] ^ m[807] ^ m[809] ^ m[812] ^ m[814] ^ m[815] ^ m[818] ^ m[819] ^ m[821] ^ m[823] ^ m[824] ^ m[827] ^ m[829] ^ m[830] ^ m[831] ^ m[834] ^ m[835] ^ m[837] ^ m[839] ^ m[841] ^ m[842] ^ m[844] ^ m[847] ^ m[848] ^ m[850] ^ m[851] ^ m[854] ^ m[855] ^ m[857] ^ m[859] ^ m[861] ^ m[862] ^ m[863] ^ m[865] ^ m[867] ^ m[869] ^ m[871] ^ m[872] ^ m[874] ^ m[877] ^ m[878] ^ m[879] ^ m[881] ^ m[883] ^ m[884] ^ m[885] ^ m[887] ^ m[889] ^ m[891] ^ m[893] ^ m[894] ^ m[896] ^ m[897] ^ m[899] ^ m[902] ^ m[903] ^ m[905] ^ m[907] ^ m[909] ^ m[911] ^ m[913] ^ m[914] ^ m[915] ^ m[917] ^ m[919] ^ m[920] ^ m[924] ^ m[925] ^ m[927] ^ m[929] ^ m[931] ^ m[932] ^ m[934] ^ m[935] ^ m[937] ^ m[940] ^ m[941] ^ m[942] ^ m[944] ^ m[946] ^ m[948] ^ m[950] ^ m[952] ^ m[954] ^ m[955] ^ m[956] ^ m[958] ^ m[959] ^ m[960] ^ m[962] ^ m[966] ^ m[967] ^ m[969] ^ m[970] ^ m[971] ^ m[973] ^ m[975] ^ m[977] ^ m[978] ^ m[979] ^ m[982] ^ m[983] ^ m[985] ^ m[987] ^ m[988] ^ m[989] ^ m[992] ^ m[993] ^ m[994] ^ m[996] ^ m[998] ^ m[999] ^ m[1001] ^ m[1002] ^ m[1003] ^ m[1005] ^ m[1007] ^ m[1008] ^ m[1009] ^ m[1010] ^ m[1012];
    assign parity[2] = m[0] ^ m[2] ^ m[4] ^ m[6] ^ m[8] ^ m[10] ^ m[12] ^ m[14] ^ m[16] ^ m[18] ^ m[20] ^ m[22] ^ m[23] ^ m[25] ^ m[28] ^ m[30] ^ m[32] ^ m[34] ^ m[36] ^ m[38] ^ m[40] ^ m[42] ^ m[44] ^ m[46] ^ m[48] ^ m[50] ^ m[51] ^ m[54] ^ m[56] ^ m[57] ^ m[60] ^ m[62] ^ m[64] ^ m[66] ^ m[68] ^ m[70] ^ m[72] ^ m[74] ^ m[75] ^ m[78] ^ m[80] ^ m[82] ^ m[84] ^ m[85] ^ m[88] ^ m[90] ^ m[92] ^ m[94] ^ m[95] ^ m[98] ^ m[100] ^ m[102] ^ m[104] ^ m[106] ^ m[108] ^ m[109] ^ m[111] ^ m[114] ^ m[116] ^ m[118] ^ m[120] ^ m[122] ^ m[123] ^ m[126] ^ m[128] ^ m[129] ^ m[132] ^ m[134] ^ m[135] ^ m[138] ^ m[139] ^ m[142] ^ m[144] ^ m[145] ^ m[148] ^ m[150] ^ m[152] ^ m[154] ^ m[156] ^ m[157] ^ m[160] ^ m[162] ^ m[163] ^ m[166] ^ m[168] ^ m[169] ^ m[172] ^ m[173] ^ m[176] ^ m[178] ^ m[180] ^ m[183] ^ m[184] ^ m[188] ^ m[192] ^ m[195] ^ m[197] ^ m[199] ^ m[202] ^ m[204] ^ m[205] ^ m[207] ^ m[211] ^ m[213] ^ m[216] ^ m[218] ^ m[221] ^ m[223] ^ m[226] ^ m[229] ^ m[231] ^ m[234] ^ m[236] ^ m[239] ^ m[240] ^ m[244] ^ m[247] ^ m[249] ^ m[250] ^ m[253] ^ m[257] ^ m[260] ^ m[261] ^ m[264] ^ m[266] ^ m[271] ^ m[273] ^ m[275] ^ m[278] ^ m[281] ^ m[282] ^ m[286] ^ m[287] ^ m[291] ^ m[292] ^ m[295] ^ m[296] ^ m[300] ^ m[301] ^ m[303] ^ m[307] ^ m[308] ^ m[311] ^ m[313] ^ m[315] ^ m[317] ^ m[318] ^ m[321] ^ m[323] ^ m[324] ^ m[327] ^ m[329] ^ m[331] ^ m[333] ^ m[335] ^ m[337] ^ m[338] ^ m[341] ^ m[343] ^ m[344] ^ m[347] ^ m[349] ^ m[351] ^ m[353] ^ m[354] ^ m[357] ^ m[359] ^ m[360] ^ m[363] ^ m[365] ^ m[366] ^ m[369] ^ m[371] ^ m[372] ^ m[375] ^ m[377] ^ m[378] ^ m[381] ^ m[382] ^ m[384] ^ m[387] ^ m[388] ^ m[391] ^ m[393] ^ m[395] ^ m[397] ^ m[399] ^ m[401] ^ m[402] ^ m[404] ^ m[407] ^ m[409] ^ m[411] ^ m[413] ^ m[415] ^ m[417] ^ m[418] ^ m[420] ^ m[423] ^ m[425] ^ m[427] ^ m[429] ^ m[430] ^ m[432] ^ m[435] ^ m[437] ^ m[439] ^ m[441] ^ m[443] ^ m[444] ^ m[446] ^ m[448] ^ m[450] ^ m[453] ^ m[455] ^ m[457] ^ m[459] ^ m[460] ^ m[462] ^ m[465] ^ m[467] ^ m[469] ^ m[470] ^ m[472] ^ m[475] ^ m[477] ^ m[479] ^ m[481] ^ m[482] ^ m[484] ^ m[487] ^ m[488] ^ m[490] ^ m[493] ^ m[495] ^ m[496] ^ m[499] ^ m[501] ^ m[502] ^ m[505] ^ m[507] ^ m[508] ^ m[511] ^ m[512] ^ m[514] ^ m[517] ^ m[519] ^ m[520] ^ m[522] ^ m[524] ^ m[526] ^ m[529] ^ m[531] ^ m[532] ^ m[535] ^ m[537] ^ m[538] ^ m[541] ^ m[542] ^ m[544] ^ m[546] ^ m[549] ^ m[550] ^ m[553] ^ m[555] ^ m[557] ^ m[558] ^ m[560] ^ m[562] ^ m[564] ^ m[565] ^ m[567] ^ m[570] ^ m[572] ^ m[574] ^ m[576] ^ m[578] ^ m[580] ^ m[582] ^ m[584] ^ m[585] ^ m[587] ^ m[590] ^ m[592] ^ m[594] ^ m[596] ^ m[597] ^ m[600] ^ m[601] ^ m[603] ^ m[606] ^ m[608] ^ m[609] ^ m[612] ^ m[614] ^ m[615] ^ m[618] ^ m[620] ^ m[621] ^ m[624] ^ m[626] ^ m[627] ^ m[630] ^ m[631] ^ m[634] ^ m[636] ^ m[637] ^ m[640] ^ m[642] ^ m[644] ^ m[646] ^ m[647] ^ m[649] ^ m[652] ^ m[653] ^ m[656] ^ m[658] ^ m[660] ^ m[662] ^ m[663] ^ m[665] ^ m[668] ^ m[670] ^ m[672] ^ m[674] ^ m[675] ^ m[677] ^ m[680] ^ m[681] ^ m[684] ^ m[686] ^ m[687] ^ m[689] ^ m[691] ^ m[693] ^ m[696] ^ m[698] ^ m[700] ^ m[701] ^ m[703] ^ m[705] ^ m[708] ^ m[710] ^ m[712] ^ m[713] ^ m[715] ^ m[718] ^ m[720] ^ m[722] ^ m[724] ^ m[725] ^ m[727] ^ m[730] ^ m[731] ^ m[734] ^ m[736] ^ m[737] ^ m[739] ^ m[741] ^ m[744] ^ m[746] ^ m[748] ^ m[749] ^ m[751] ^ m[754] ^ m[755] ^ m[758] ^ m[760] ^ m[761] ^ m[763] ^ m[765] ^ m[767] ^ m[770] ^ m[772] ^ m[773] ^ m[775] ^ m[777] ^ m[780] ^ m[782] ^ m[784] ^ m[785] ^ m[787] ^ m[789] ^ m[792] ^ m[794] ^ m[796] ^ m[798] ^ m[799] ^ m[801] ^ m[803] ^ m[805] ^ m[808] ^ m[810] ^ m[812] ^ m[813] ^ m[815] ^ m[818] ^ m[819] ^ m[820] ^ m[822] ^ m[825] ^ m[827] ^ m[828] ^ m[830] ^ m[832] ^ m[833] ^ m[835] ^ m[837] ^ m[838] ^ m[841] ^ m[843] ^ m[845] ^ m[847] ^ m[848] ^ m[850] ^ m[852] ^ m[853] ^ m[854] ^ m[857] ^ m[858] ^ m[861] ^ m[862] ^ m[864] ^ m[865] ^ m[866] ^ m[868] ^ m[871] ^ m[873] ^ m[875] ^ m[876] ^ m[878] ^ m[879] ^ m[880] ^ m[882] ^ m[885] ^ m[886] ^ m[888] ^ m[890] ^ m[891] ^ m[892] ^ m[894] ^ m[896] ^ m[898] ^ m[899] ^ m[902] ^ m[903] ^ m[904] ^ m[907] ^ m[908] ^ m[911] ^ m[912] ^ m[914] ^ m[916] ^ m[918] ^ m[919] ^ m[921] ^ m[923] ^ m[926] ^ m[927] ^ m[929] ^ m[930] ^ m[932] ^ m[933] ^ m[935] ^ m[938] ^ m[939] ^ m[941] ^ m[942] ^ m[944] ^ m[947] ^ m[949] ^ m[950] ^ m[952] ^ m[953] ^ m[956] ^ m[957] ^ m[958] ^ m[959] ^ m[960] ^ m[963] ^ m[965] ^ m[967] ^ m[968] ^ m[970] ^ m[972] ^ m[973] ^ m[974] ^ m[977] ^ m[978] ^ m[980] ^ m[981] ^ m[982] ^ m[985] ^ m[986] ^ m[989] ^ m[990] ^ m[992] ^ m[994] ^ m[995] ^ m[997] ^ m[998] ^ m[999] ^ m[1000] ^ m[1002] ^ m[1004] ^ m[1005] ^ m[1006] ^ m[1007] ^ m[1009] ^ m[1010] ^ m[1011];
    assign parity[3] = m[0] ^ m[2] ^ m[4] ^ m[6] ^ m[8] ^ m[10] ^ m[12] ^ m[14] ^ m[16] ^ m[18] ^ m[19] ^ m[21] ^ m[24] ^ m[26] ^ m[28] ^ m[30] ^ m[32] ^ m[34] ^ m[36] ^ m[38] ^ m[40] ^ m[42] ^ m[44] ^ m[46] ^ m[47] ^ m[50] ^ m[52] ^ m[53] ^ m[56] ^ m[58] ^ m[60] ^ m[62] ^ m[64] ^ m[66] ^ m[68] ^ m[70] ^ m[71] ^ m[74] ^ m[76] ^ m[78] ^ m[80] ^ m[81] ^ m[84] ^ m[86] ^ m[88] ^ m[90] ^ m[91] ^ m[94] ^ m[96] ^ m[98] ^ m[100] ^ m[102] ^ m[104] ^ m[105] ^ m[107] ^ m[110] ^ m[112] ^ m[114] ^ m[116] ^ m[118] ^ m[120] ^ m[122] ^ m[123] ^ m[125] ^ m[127] ^ m[130] ^ m[131] ^ m[134] ^ m[136] ^ m[138] ^ m[140] ^ m[141] ^ m[144] ^ m[146] ^ m[148] ^ m[150] ^ m[152] ^ m[154] ^ m[156] ^ m[157] ^ m[159] ^ m[161] ^ m[164] ^ m[165] ^ m[168] ^ m[170] ^ m[172] ^ m[174] ^ m[176] ^ m[178] ^ m[180] ^ m[181] ^ m[185] ^ m[189] ^ m[192] ^ m[194] ^ m[197] ^ m[199] ^ m[200] ^ m[204] ^ m[206] ^ m[209] ^ m[210] ^ m[213] ^ m[215] ^ m[219] ^ m[220] ^ m[224] ^ m[227] ^ m[229] ^ m[231] ^ m[233] ^ m[236] ^ m[239] ^ m[240] ^ m[243] ^ m[247] ^ m[248] ^ m[251] ^ m[255] ^ m[258] ^ m[259] ^ m[262] ^ m[264] ^ m[266] ^ m[269] ^ m[272] ^ m[276] ^ m[277] ^ m[280] ^ m[283] ^ m[286] ^ m[289] ^ m[290] ^ m[294] ^ m[295] ^ m[297] ^ m[300] ^ m[301] ^ m[303] ^ m[306] ^ m[309] ^ m[311] ^ m[313] ^ m[314] ^ m[317] ^ m[319] ^ m[320] ^ m[323] ^ m[325] ^ m[327] ^ m[329] ^ m[331] ^ m[333] ^ m[334] ^ m[337] ^ m[339] ^ m[340] ^ m[343] ^ m[345] ^ m[347] ^ m[349] ^ m[350] ^ m[353] ^ m[355] ^ m[356] ^ m[359] ^ m[361] ^ m[363] ^ m[365] ^ m[366] ^ m[369] ^ m[370] ^ m[372] ^ m[374] ^ m[376] ^ m[379] ^ m[380] ^ m[383] ^ m[385] ^ m[387] ^ m[389] ^ m[391] ^ m[393] ^ m[395] ^ m[397] ^ m[398] ^ m[400] ^ m[403] ^ m[405] ^ m[407] ^ m[409] ^ m[411] ^ m[413] ^ m[415] ^ m[416] ^ m[419] ^ m[421] ^ m[423] ^ m[425] ^ m[426] ^ m[429] ^ m[431] ^ m[432] ^ m[435] ^ m[436] ^ m[438] ^ m[440] ^ m[442] ^ m[445] ^ m[447] ^ m[449] ^ m[451] ^ m[453] ^ m[455] ^ m[456] ^ m[458] ^ m[461] ^ m[463] ^ m[465] ^ m[466] ^ m[469] ^ m[471] ^ m[472] ^ m[475] ^ m[476] ^ m[479] ^ m[480] ^ m[482] ^ m[485] ^ m[486] ^ m[489] ^ m[491] ^ m[493] ^ m[495] ^ m[496] ^ m[498] ^ m[500] ^ m[503] ^ m[504] ^ m[507] ^ m[509] ^ m[511] ^ m[513] ^ m[514] ^ m[517] ^ m[518] ^ m[520] ^ m[523] ^ m[524] ^ m[527] ^ m[528] ^ m[531] ^ m[533] ^ m[534] ^ m[537] ^ m[539] ^ m[540] ^ m[543] ^ m[545] ^ m[546] ^ m[549] ^ m[550] ^ m[553] ^ m[554] ^ m[557] ^ m[558] ^ m[560] ^ m[561] ^ m[563] ^ m[566] ^ m[568] ^ m[570] ^ m[572] ^ m[574] ^ m[576] ^ m[577] ^ m[580] ^ m[582] ^ m[583] ^ m[585] ^ m[588] ^ m[589] ^ m[592] ^ m[593] ^ m[596] ^ m[598] ^ m[599] ^ m[602] ^ m[604] ^ m[606] ^ m[608] ^ m[610] ^ m[612] ^ m[614] ^ m[615] ^ m[617] ^ m[619] ^ m[622] ^ m[623] ^ m[626] ^ m[628] ^ m[630] ^ m[632] ^ m[634] ^ m[636] ^ m[637] ^ m[640] ^ m[641] ^ m[643] ^ m[645] ^ m[648] ^ m[650] ^ m[652] ^ m[654] ^ m[656] ^ m[657] ^ m[659] ^ m[662] ^ m[664] ^ m[665] ^ m[668] ^ m[669] ^ m[672] ^ m[673] ^ m[675] ^ m[678] ^ m[679] ^ m[682] ^ m[683] ^ m[686] ^ m[688] ^ m[689] ^ m[692] ^ m[693] ^ m[696] ^ m[697] ^ m[699] ^ m[702] ^ m[704] ^ m[706] ^ m[708] ^ m[709] ^ m[712] ^ m[714] ^ m[715] ^ m[718] ^ m[719] ^ m[722] ^ m[723] ^ m[725] ^ m[728] ^ m[729] ^ m[732] ^ m[733] ^ m[736] ^ m[738] ^ m[739] ^ m[742] ^ m[743] ^ m[746] ^ m[747] ^ m[749] ^ m[752] ^ m[753] ^ m[756] ^ m[757] ^ m[760] ^ m[762] ^ m[763] ^ m[766] ^ m[767] ^ m[770] ^ m[771] ^ m[773] ^ m[776] ^ m[777] ^ m[780] ^ m[781] ^ m[784] ^ m[786] ^ m[787] ^ m[789] ^ m[791] ^ m[793] ^ m[795] ^ m[797] ^ m[800] ^ m[802] ^ m[804] ^ m[806] ^ m[808] ^ m[810] ^ m[811] ^ m[813] ^ m[815] ^ m[817] ^ m[819] ^ m[821] ^ m[822] ^ m[825] ^ m[827] ^ m[829] ^ m[830] ^ m[831] ^ m[833] ^ m[835] ^ m[837] ^ m[838] ^ m[840] ^ m[843] ^ m[844] ^ m[846] ^ m[848] ^ m[850] ^ m[851] ^ m[853] ^ m[855] ^ m[856] ^ m[858] ^ m[860] ^ m[862] ^ m[863] ^ m[865] ^ m[867] ^ m[869] ^ m[870] ^ m[873] ^ m[875] ^ m[876] ^ m[877] ^ m[880] ^ m[881] ^ m[883] ^ m[885] ^ m[886] ^ m[888] ^ m[889] ^ m[890] ^ m[892] ^ m[893] ^ m[896] ^ m[897] ^ m[900] ^ m[902] ^ m[903] ^ m[905] ^ m[906] ^ m[909] ^ m[910] ^ m[912] ^ m[914] ^ m[916] ^ m[917] ^ m[918] ^ m[922] ^ m[923] ^ m[925] ^ m[927] ^ m[928] ^ m[930] ^ m[932] ^ m[934] ^ m[936] ^ m[938] ^ m[939] ^ m[940] ^ m[943] ^ m[944] ^ m[946] ^ m[947] ^ m[949] ^ m[951] ^ m[952] ^ m[954] ^ m[955] ^ m[959] ^ m[960] ^ m[961] ^ m[962] ^ m[964] ^ m[967] ^ m[968] ^ m[970] ^ m[971] ^ m[972] ^ m[974] ^ m[976] ^ m[978] ^ m[980] ^ m[982] ^ m[983] ^ m[984] ^ m[987] ^ m[989] ^ m[990] ^ m[991] ^ m[994] ^ m[995] ^ m[997] ^ m[998] ^ m[999] ^ m[1000] ^ m[1001] ^ m[1003] ^ m[1004] ^ m[1007] ^ m[1008] ^ m[1010] ^ m[1011] ^ m[1012];
    assign parity[4] = m[0] ^ m[2] ^ m[4] ^ m[6] ^ m[8] ^ m[10] ^ m[12] ^ m[14] ^ m[15] ^ m[17] ^ m[20] ^ m[22] ^ m[24] ^ m[26] ^ m[28] ^ m[30] ^ m[32] ^ m[34] ^ m[36] ^ m[38] ^ m[40] ^ m[42] ^ m[43] ^ m[46] ^ m[48] ^ m[49] ^ m[52] ^ m[54] ^ m[56] ^ m[58] ^ m[60] ^ m[62] ^ m[64] ^ m[66] ^ m[67] ^ m[70] ^ m[72] ^ m[74] ^ m[76] ^ m[77] ^ m[80] ^ m[82] ^ m[84] ^ m[86] ^ m[87] ^ m[90] ^ m[92] ^ m[94] ^ m[96] ^ m[98] ^ m[100] ^ m[101] ^ m[104] ^ m[106] ^ m[107] ^ m[110] ^ m[111] ^ m[114] ^ m[115] ^ m[118] ^ m[119] ^ m[121] ^ m[124] ^ m[126] ^ m[128] ^ m[130] ^ m[132] ^ m[134] ^ m[136] ^ m[138] ^ m[140] ^ m[141] ^ m[144] ^ m[145] ^ m[148] ^ m[149] ^ m[152] ^ m[153] ^ m[155] ^ m[158] ^ m[160] ^ m[162] ^ m[164] ^ m[166] ^ m[168] ^ m[170] ^ m[172] ^ m[174] ^ m[176] ^ m[178] ^ m[179] ^ m[182] ^ m[186] ^ m[189] ^ m[192] ^ m[193] ^ m[196] ^ m[199] ^ m[201] ^ m[204] ^ m[206] ^ m[209] ^ m[211] ^ m[213] ^ m[215] ^ m[218] ^ m[220] ^ m[223] ^ m[227] ^ m[228] ^ m[230] ^ m[232] ^ m[235] ^ m[237] ^ m[242] ^ m[245] ^ m[247] ^ m[249] ^ m[251] ^ m[254] ^ m[257] ^ m[259] ^ m[261] ^ m[263] ^ m[267] ^ m[270] ^ m[274] ^ m[277] ^ m[279] ^ m[281] ^ m[283] ^ m[286] ^ m[289] ^ m[290] ^ m[292] ^ m[295] ^ m[296] ^ m[299] ^ m[302] ^ m[305] ^ m[307] ^ m[309] ^ m[310] ^ m[313] ^ m[315] ^ m[316] ^ m[319] ^ m[321] ^ m[323] ^ m[325] ^ m[327] ^ m[329] ^ m[330] ^ m[333] ^ m[335] ^ m[336] ^ m[339] ^ m[341] ^ m[343] ^ m[345] ^ m[347] ^ m[349] ^ m[350] ^ m[353] ^ m[354] ^ m[356] ^ m[358] ^ m[360] ^ m[362] ^ m[364] ^ m[367] ^ m[368] ^ m[371] ^ m[373] ^ m[375] ^ m[377] ^ m[379] ^ m[381] ^ m[383] ^ m[385] ^ m[387] ^ m[389] ^ m[391] ^ m[393] ^ m[394] ^ m[396] ^ m[399] ^ m[401] ^ m[403] ^ m[405] ^ m[407] ^ m[409] ^ m[411] ^ m[413] ^ m[414] ^ m[416] ^ m[419] ^ m[420] ^ m[423] ^ m[424] ^ m[426] ^ m[428] ^ m[430] ^ m[433] ^ m[434] ^ m[437] ^ m[439] ^ m[441] ^ m[443] ^ m[445] ^ m[447] ^ m[449] ^ m[451] ^ m[453] ^ m[455] ^ m[456] ^ m[459] ^ m[460] ^ m[463] ^ m[464] ^ m[466] ^ m[468] ^ m[470] ^ m[473] ^ m[474] ^ m[477] ^ m[478] ^ m[481] ^ m[483] ^ m[485] ^ m[487] ^ m[489] ^ m[491] ^ m[493] ^ m[495] ^ m[496] ^ m[498] ^ m[500] ^ m[502] ^ m[504] ^ m[506] ^ m[508] ^ m[510] ^ m[512] ^ m[515] ^ m[516] ^ m[519] ^ m[521] ^ m[523] ^ m[525] ^ m[527] ^ m[529] ^ m[531] ^ m[533] ^ m[534] ^ m[536] ^ m[538] ^ m[541] ^ m[542] ^ m[545] ^ m[547] ^ m[549] ^ m[551] ^ m[553] ^ m[555] ^ m[557] ^ m[558] ^ m[559] ^ m[561] ^ m[564] ^ m[565] ^ m[568] ^ m[569] ^ m[572] ^ m[573] ^ m[576] ^ m[578] ^ m[579] ^ m[581] ^ m[584] ^ m[586] ^ m[588] ^ m[590] ^ m[592] ^ m[594] ^ m[596] ^ m[598] ^ m[599] ^ m[602] ^ m[603] ^ m[606] ^ m[607] ^ m[610] ^ m[611] ^ m[614] ^ m[616] ^ m[617] ^ m[620] ^ m[621] ^ m[624] ^ m[626] ^ m[628] ^ m[629] ^ m[632] ^ m[633] ^ m[636] ^ m[638] ^ m[639] ^ m[642] ^ m[644] ^ m[646] ^ m[648] ^ m[650] ^ m[652] ^ m[654] ^ m[656] ^ m[657] ^ m[659] ^ m[662] ^ m[663] ^ m[665] ^ m[667] ^ m[669] ^ m[671] ^ m[673] ^ m[676] ^ m[677] ^ m[680] ^ m[681] ^ m[684] ^ m[685] ^ m[688] ^ m[690] ^ m[692] ^ m[694] ^ m[696] ^ m[698] ^ m[699] ^ m[701] ^ m[703] ^ m[706] ^ m[707] ^ m[709] ^ m[711] ^ m[713] ^ m[716] ^ m[717] ^ m[720] ^ m[721] ^ m[724] ^ m[726] ^ m[728] ^ m[730] ^ m[732] ^ m[734] ^ m[736] ^ m[738] ^ m[739] ^ m[742] ^ m[743] ^ m[746] ^ m[747] ^ m[749] ^ m[751] ^ m[753] ^ m[755] ^ m[757] ^ m[759] ^ m[761] ^ m[764] ^ m[765] ^ m[768] ^ m[769] ^ m[772] ^ m[774] ^ m[776] ^ m[778] ^ m[779] ^ m[782] ^ m[783] ^ m[786] ^ m[788] ^ m[789] ^ m[792] ^ m[793] ^ m[796] ^ m[797] ^ m[800] ^ m[801] ^ m[804] ^ m[805] ^ m[808] ^ m[809] ^ m[811] ^ m[813] ^ m[816] ^ m[817] ^ m[819] ^ m[820] ^ m[823] ^ m[824] ^ m[826] ^ m[828] ^ m[830] ^ m[831] ^ m[833] ^ m[835] ^ m[836] ^ m[839] ^ m[841] ^ m[842] ^ m[845] ^ m[847] ^ m[848] ^ m[849] ^ m[851] ^ m[853] ^ m[855] ^ m[856] ^ m[859] ^ m[860] ^ m[861] ^ m[864] ^ m[865] ^ m[866] ^ m[869] ^ m[871] ^ m[872] ^ m[875] ^ m[876] ^ m[878] ^ m[880] ^ m[881] ^ m[883] ^ m[884] ^ m[886] ^ m[888] ^ m[890] ^ m[891] ^ m[893] ^ m[894] ^ m[895] ^ m[897] ^ m[900] ^ m[902] ^ m[904] ^ m[905] ^ m[906] ^ m[908] ^ m[910] ^ m[911] ^ m[914] ^ m[915] ^ m[918] ^ m[920] ^ m[921] ^ m[923] ^ m[925] ^ m[926] ^ m[928] ^ m[929] ^ m[931] ^ m[933] ^ m[935] ^ m[937] ^ m[939] ^ m[941] ^ m[943] ^ m[945] ^ m[947] ^ m[948] ^ m[950] ^ m[952] ^ m[953] ^ m[955] ^ m[956] ^ m[958] ^ m[959] ^ m[961] ^ m[962] ^ m[964] ^ m[965] ^ m[969] ^ m[970] ^ m[971] ^ m[973] ^ m[975] ^ m[976] ^ m[978] ^ m[979] ^ m[980] ^ m[981] ^ m[985] ^ m[986] ^ m[987] ^ m[989] ^ m[991] ^ m[993] ^ m[995] ^ m[997] ^ m[998] ^ m[1000] ^ m[1001] ^ m[1002] ^ m[1003] ^ m[1004] ^ m[1006] ^ m[1007] ^ m[1008] ^ m[1009] ^ m[1011];
    assign parity[5] = m[0] ^ m[2] ^ m[4] ^ m[6] ^ m[8] ^ m[10] ^ m[11] ^ m[13] ^ m[16] ^ m[18] ^ m[20] ^ m[22] ^ m[24] ^ m[26] ^ m[28] ^ m[30] ^ m[32] ^ m[34] ^ m[36] ^ m[38] ^ m[39] ^ m[42] ^ m[44] ^ m[45] ^ m[48] ^ m[50] ^ m[52] ^ m[54] ^ m[56] ^ m[58] ^ m[60] ^ m[62] ^ m[63] ^ m[66] ^ m[68] ^ m[70] ^ m[72] ^ m[73] ^ m[76] ^ m[78] ^ m[80] ^ m[82] ^ m[84] ^ m[86] ^ m[87] ^ m[90] ^ m[91] ^ m[94] ^ m[95] ^ m[97] ^ m[99] ^ m[102] ^ m[103] ^ m[106] ^ m[108] ^ m[110] ^ m[112] ^ m[114] ^ m[116] ^ m[118] ^ m[120] ^ m[121] ^ m[124] ^ m[125] ^ m[128] ^ m[129] ^ m[132] ^ m[133] ^ m[136] ^ m[137] ^ m[140] ^ m[142] ^ m[144] ^ m[146] ^ m[148] ^ m[150] ^ m[151] ^ m[154] ^ m[156] ^ m[158] ^ m[160] ^ m[162] ^ m[164] ^ m[166] ^ m[168] ^ m[170] ^ m[172] ^ m[174] ^ m[175] ^ m[178] ^ m[180] ^ m[182] ^ m[185] ^ m[188] ^ m[191] ^ m[193] ^ m[196] ^ m[198] ^ m[200] ^ m[203] ^ m[206] ^ m[207] ^ m[210] ^ m[213] ^ m[214] ^ m[217] ^ m[222] ^ m[225] ^ m[226] ^ m[229] ^ m[232] ^ m[234] ^ m[236] ^ m[238] ^ m[242] ^ m[245] ^ m[246] ^ m[249] ^ m[252] ^ m[255] ^ m[258] ^ m[259] ^ m[261] ^ m[264] ^ m[267] ^ m[270] ^ m[273] ^ m[276] ^ m[278] ^ m[280] ^ m[284] ^ m[287] ^ m[288] ^ m[289] ^ m[294] ^ m[295] ^ m[298] ^ m[300] ^ m[302] ^ m[304] ^ m[307] ^ m[309] ^ m[311] ^ m[312] ^ m[315] ^ m[317] ^ m[319] ^ m[321] ^ m[323] ^ m[325] ^ m[327] ^ m[329] ^ m[330] ^ m[333] ^ m[334] ^ m[336] ^ m[338] ^ m[340] ^ m[342] ^ m[344] ^ m[346] ^ m[348] ^ m[351] ^ m[352] ^ m[355] ^ m[357] ^ m[359] ^ m[361] ^ m[363] ^ m[365] ^ m[367] ^ m[369] ^ m[371] ^ m[373] ^ m[375] ^ m[377] ^ m[379] ^ m[381] ^ m[383] ^ m[385] ^ m[387] ^ m[389] ^ m[390] ^ m[393] ^ m[395] ^ m[396] ^ m[399] ^ m[400] ^ m[403] ^ m[404] ^ m[407] ^ m[408] ^ m[411] ^ m[412] ^ m[414] ^ m[417] ^ m[418] ^ m[421] ^ m[422] ^ m[425] ^ m[427] ^ m[429] ^ m[431] ^ m[433] ^ m[435] ^ m[437] ^ m[439] ^ m[441] ^ m[443] ^ m[445] ^ m[447] ^ m[449] ^ m[451] ^ m[453] ^ m[455] ^ m[456] ^ m[458] ^ m[460] ^ m[462] ^ m[464] ^ m[467] ^ m[468] ^ m[471] ^ m[472] ^ m[475] ^ m[476] ^ m[479] ^ m[480] ^ m[483] ^ m[484] ^ m[487] ^ m[488] ^ m[491] ^ m[492] ^ m[495] ^ m[497] ^ m[498] ^ m[501] ^ m[502] ^ m[505] ^ m[506] ^ m[509] ^ m[510] ^ m[513] ^ m[514] ^ m[517] ^ m[518] ^ m[521] ^ m[522] ^ m[525] ^ m[526] ^ m[529] ^ m[530] ^ m[533] ^ m[535] ^ m[536] ^ m[539] ^ m[540] ^ m[543] ^ m[544] ^ m[547] ^ m[548] ^ m[551] ^ m[552] ^ m[555] ^ m[556] ^ m[558] ^ m[560] ^ m[562] ^ m[564] ^ m[566] ^ m[568] ^ m[569] ^ m[572] ^ m[574] ^ m[576] ^ m[577] ^ m[579] ^ m[582] ^ m[583] ^ m[586] ^ m[587] ^ m[590] ^ m[591] ^ m[594] ^ m[595] ^ m[598] ^ m[600] ^ m[602] ^ m[604] ^ m[606] ^ m[608] ^ m[609] ^ m[612] ^ m[613] ^ m[616] ^ m[617] ^ m[620] ^ m[621] ^ m[624] ^ m[625] ^ m[628] ^ m[629] ^ m[632] ^ m[633] ^ m[636] ^ m[637] ^ m[639] ^ m[641] ^ m[643] ^ m[645] ^ m[647] ^ m[649] ^ m[651] ^ m[653] ^ m[655] ^ m[658] ^ m[660] ^ m[661] ^ m[664] ^ m[666] ^ m[668] ^ m[670] ^ m[672] ^ m[674] ^ m[676] ^ m[678] ^ m[680] ^ m[682] ^ m[684] ^ m[686] ^ m[688] ^ m[690] ^ m[692] ^ m[694] ^ m[696] ^ m[698] ^ m[699] ^ m[702] ^ m[703] ^ m[706] ^ m[707] ^ m[709] ^ m[711] ^ m[713] ^ m[715] ^ m[717] ^ m[719] ^ m[721] ^ m[723] ^ m[725] ^ m[727] ^ m[729] ^ m[731] ^ m[733] ^ m[735] ^ m[737] ^ m[740] ^ m[741] ^ m[744] ^ m[745] ^ m[748] ^ m[750] ^ m[752] ^ m[754] ^ m[756] ^ m[758] ^ m[760] ^ m[762] ^ m[764] ^ m[766] ^ m[768] ^ m[770] ^ m[772] ^ m[774] ^ m[776] ^ m[778] ^ m[780] ^ m[782] ^ m[784] ^ m[786] ^ m[788] ^ m[789] ^ m[792] ^ m[793] ^ m[796] ^ m[797] ^ m[800] ^ m[801] ^ m[804] ^ m[805] ^ m[808] ^ m[809] ^ m[811] ^ m[812] ^ m[815] ^ m[817] ^ m[818] ^ m[820] ^ m[822] ^ m[824] ^ m[826] ^ m[828] ^ m[829] ^ m[830] ^ m[833] ^ m[834] ^ m[836] ^ m[838] ^ m[840] ^ m[842] ^ m[844] ^ m[845] ^ m[846] ^ m[849] ^ m[851] ^ m[852] ^ m[854] ^ m[857] ^ m[858] ^ m[860] ^ m[862] ^ m[863] ^ m[865] ^ m[867] ^ m[868] ^ m[870] ^ m[873] ^ m[874] ^ m[876] ^ m[878] ^ m[879] ^ m[880] ^ m[882] ^ m[884] ^ m[886] ^ m[887] ^ m[889] ^ m[891] ^ m[893] ^ m[895] ^ m[896] ^ m[898] ^ m[900] ^ m[901] ^ m[904] ^ m[905] ^ m[907] ^ m[909] ^ m[911] ^ m[913] ^ m[914] ^ m[916] ^ m[918] ^ m[920] ^ m[922] ^ m[923] ^ m[924] ^ m[925] ^ m[928] ^ m[930] ^ m[931] ^ m[933] ^ m[935] ^ m[937] ^ m[938] ^ m[940] ^ m[942] ^ m[944] ^ m[946] ^ m[949] ^ m[950] ^ m[951] ^ m[953] ^ m[956] ^ m[957] ^ m[959] ^ m[961] ^ m[963] ^ m[964] ^ m[966] ^ m[967] ^ m[969] ^ m[970] ^ m[971] ^ m[972] ^ m[975] ^ m[976] ^ m[977] ^ m[979] ^ m[981] ^ m[983] ^ m[984] ^ m[986] ^ m[988] ^ m[990] ^ m[992] ^ m[993] ^ m[995] ^ m[996] ^ m[998] ^ m[999] ^ m[1001] ^ m[1002] ^ m[1003] ^ m[1005] ^ m[1006] ^ m[1008] ^ m[1010] ^ m[1011] ^ m[1012];
    assign parity[6] = m[0] ^ m[2] ^ m[4] ^ m[6] ^ m[7] ^ m[9] ^ m[12] ^ m[14] ^ m[16] ^ m[18] ^ m[20] ^ m[22] ^ m[24] ^ m[26] ^ m[28] ^ m[30] ^ m[32] ^ m[34] ^ m[35] ^ m[38] ^ m[40] ^ m[41] ^ m[44] ^ m[46] ^ m[48] ^ m[50] ^ m[52] ^ m[54] ^ m[56] ^ m[58] ^ m[60] ^ m[62] ^ m[63] ^ m[66] ^ m[67] ^ m[69] ^ m[71] ^ m[74] ^ m[75] ^ m[78] ^ m[79] ^ m[82] ^ m[83] ^ m[86] ^ m[88] ^ m[90] ^ m[92] ^ m[94] ^ m[96] ^ m[97] ^ m[100] ^ m[101] ^ m[104] ^ m[105] ^ m[108] ^ m[109] ^ m[112] ^ m[113] ^ m[116] ^ m[117] ^ m[120] ^ m[122] ^ m[124] ^ m[126] ^ m[128] ^ m[130] ^ m[132] ^ m[134] ^ m[136] ^ m[138] ^ m[140] ^ m[142] ^ m[144] ^ m[146] ^ m[147] ^ m[150] ^ m[152] ^ m[154] ^ m[156] ^ m[158] ^ m[160] ^ m[162] ^ m[164] ^ m[166] ^ m[168] ^ m[170] ^ m[172] ^ m[174] ^ m[175] ^ m[178] ^ m[179] ^ m[181] ^ m[184] ^ m[187] ^ m[190] ^ m[194] ^ m[196] ^ m[198] ^ m[201] ^ m[202] ^ m[205] ^ m[208] ^ m[210] ^ m[212] ^ m[216] ^ m[219] ^ m[222] ^ m[225] ^ m[226] ^ m[229] ^ m[232] ^ m[234] ^ m[236] ^ m[238] ^ m[242] ^ m[245] ^ m[246] ^ m[249] ^ m[251] ^ m[254] ^ m[257] ^ m[258] ^ m[260] ^ m[263] ^ m[266] ^ m[269] ^ m[272] ^ m[275] ^ m[277] ^ m[279] ^ m[282] ^ m[285] ^ m[287] ^ m[291] ^ m[293] ^ m[295] ^ m[298] ^ m[300] ^ m[302] ^ m[304] ^ m[307] ^ m[309] ^ m[310] ^ m[312] ^ m[314] ^ m[316] ^ m[318] ^ m[320] ^ m[322] ^ m[324] ^ m[326] ^ m[328] ^ m[331] ^ m[332] ^ m[335] ^ m[337] ^ m[339] ^ m[341] ^ m[343] ^ m[345] ^ m[347] ^ m[349] ^ m[351] ^ m[353] ^ m[355] ^ m[357] ^ m[359] ^ m[361] ^ m[363] ^ m[365] ^ m[367] ^ m[369] ^ m[371] ^ m[373] ^ m[375] ^ m[377] ^ m[379] ^ m[381] ^ m[383] ^ m[385] ^ m[387] ^ m[389] ^ m[390] ^ m[393] ^ m[394] ^ m[396] ^ m[398] ^ m[400] ^ m[402] ^ m[404] ^ m[406] ^ m[408] ^ m[410] ^ m[412] ^ m[415] ^ m[416] ^ m[419] ^ m[420] ^ m[423] ^ m[424] ^ m[427] ^ m[428] ^ m[431] ^ m[432] ^ m[435] ^ m[436] ^ m[439] ^ m[440] ^ m[443] ^ m[444] ^ m[447] ^ m[448] ^ m[451] ^ m[452] ^ m[455] ^ m[457] ^ m[458] ^ m[461] ^ m[462] ^ m[465] ^ m[466] ^ m[469] ^ m[470] ^ m[473] ^ m[474] ^ m[477] ^ m[478] ^ m[481] ^ m[482] ^ m[485] ^ m[486] ^ m[489] ^ m[490] ^ m[493] ^ m[494] ^ m[497] ^ m[499] ^ m[501] ^ m[503] ^ m[505] ^ m[507] ^ m[509] ^ m[511] ^ m[513] ^ m[515] ^ m[517] ^ m[519] ^ m[521] ^ m[523] ^ m[525] ^ m[527] ^ m[529] ^ m[531] ^ m[533] ^ m[535] ^ m[536] ^ m[539] ^ m[540] ^ m[543] ^ m[544] ^ m[547] ^ m[548] ^ m[551] ^ m[552] ^ m[555] ^ m[556] ^ m[558] ^ m[559] ^ m[561] ^ m[563] ^ m[565] ^ m[567] ^ m[569] ^ m[571] ^ m[573] ^ m[575] ^ m[577] ^ m[580] ^ m[581] ^ m[584] ^ m[585] ^ m[588] ^ m[589] ^ m[592] ^ m[593] ^ m[596] ^ m[597] ^ m[600] ^ m[601] ^ m[604] ^ m[605] ^ m[608] ^ m[609] ^ m[612] ^ m[613] ^ m[616] ^ m[618] ^ m[620] ^ m[622] ^ m[624] ^ m[625] ^ m[628] ^ m[630] ^ m[632] ^ m[634] ^ m[636] ^ m[638] ^ m[639] ^ m[642] ^ m[643] ^ m[646] ^ m[647] ^ m[650] ^ m[651] ^ m[654] ^ m[655] ^ m[657] ^ m[659] ^ m[662] ^ m[663] ^ m[666] ^ m[667] ^ m[670] ^ m[671] ^ m[674] ^ m[675] ^ m[678] ^ m[679] ^ m[682] ^ m[683] ^ m[686] ^ m[687] ^ m[690] ^ m[691] ^ m[694] ^ m[695] ^ m[698] ^ m[700] ^ m[701] ^ m[704] ^ m[706] ^ m[708] ^ m[709] ^ m[712] ^ m[713] ^ m[716] ^ m[717] ^ m[720] ^ m[721] ^ m[724] ^ m[725] ^ m[728] ^ m[729] ^ m[732] ^ m[733] ^ m[736] ^ m[737] ^ m[740] ^ m[741] ^ m[744] ^ m[745] ^ m[748] ^ m[749] ^ m[752] ^ m[753] ^ m[756] ^ m[757] ^ m[760] ^ m[761] ^ m[764] ^ m[765] ^ m[768] ^ m[769] ^ m[772] ^ m[773] ^ m[776] ^ m[777] ^ m[779] ^ m[781] ^ m[783] ^ m[785] ^ m[787] ^ m[790] ^ m[791] ^ m[794] ^ m[795] ^ m[798] ^ m[799] ^ m[802] ^ m[803] ^ m[806] ^ m[807] ^ m[810] ^ m[812] ^ m[814] ^ m[816] ^ m[817] ^ m[819] ^ m[821] ^ m[823] ^ m[825] ^ m[826] ^ m[828] ^ m[830] ^ m[832] ^ m[833] ^ m[835] ^ m[837] ^ m[839] ^ m[840] ^ m[842] ^ m[845] ^ m[847] ^ m[848] ^ m[849] ^ m[851] ^ m[853] ^ m[855] ^ m[857] ^ m[858] ^ m[860] ^ m[862] ^ m[863] ^ m[864] ^ m[867] ^ m[868] ^ m[870] ^ m[873] ^ m[874] ^ m[876] ^ m[878] ^ m[879] ^ m[881] ^ m[882] ^ m[884] ^ m[886] ^ m[887] ^ m[889] ^ m[890] ^ m[893] ^ m[894] ^ m[897] ^ m[898] ^ m[900] ^ m[901] ^ m[903] ^ m[905] ^ m[906] ^ m[908] ^ m[910] ^ m[912] ^ m[913] ^ m[915] ^ m[917] ^ m[919] ^ m[921] ^ m[924] ^ m[926] ^ m[927] ^ m[929] ^ m[930] ^ m[932] ^ m[934] ^ m[936] ^ m[937] ^ m[939] ^ m[941] ^ m[943] ^ m[945] ^ m[946] ^ m[948] ^ m[950] ^ m[951] ^ m[954] ^ m[956] ^ m[957] ^ m[959] ^ m[961] ^ m[962] ^ m[964] ^ m[965] ^ m[967] ^ m[968] ^ m[969] ^ m[972] ^ m[973] ^ m[974] ^ m[975] ^ m[978] ^ m[980] ^ m[981] ^ m[983] ^ m[984] ^ m[985] ^ m[986] ^ m[987] ^ m[988] ^ m[990] ^ m[991] ^ m[992] ^ m[993] ^ m[994] ^ m[996] ^ m[998] ^ m[1000] ^ m[1001] ^ m[1005] ^ m[1007] ^ m[1009] ^ m[1010] ^ m[1011];
    assign parity[7] = m[0] ^ m[2] ^ m[3] ^ m[5] ^ m[8] ^ m[10] ^ m[12] ^ m[14] ^ m[16] ^ m[18] ^ m[20] ^ m[22] ^ m[24] ^ m[26] ^ m[28] ^ m[30] ^ m[32] ^ m[34] ^ m[35] ^ m[37] ^ m[39] ^ m[42] ^ m[43] ^ m[46] ^ m[47] ^ m[50] ^ m[51] ^ m[54] ^ m[55] ^ m[58] ^ m[59] ^ m[62] ^ m[64] ^ m[66] ^ m[68] ^ m[69] ^ m[72] ^ m[73] ^ m[76] ^ m[77] ^ m[80] ^ m[81] ^ m[84] ^ m[85] ^ m[88] ^ m[89] ^ m[92] ^ m[93] ^ m[96] ^ m[98] ^ m[100] ^ m[102] ^ m[104] ^ m[106] ^ m[108] ^ m[110] ^ m[112] ^ m[114] ^ m[116] ^ m[118] ^ m[120] ^ m[122] ^ m[124] ^ m[126] ^ m[128] ^ m[130] ^ m[132] ^ m[134] ^ m[136] ^ m[138] ^ m[140] ^ m[142] ^ m[144] ^ m[146] ^ m[147] ^ m[150] ^ m[151] ^ m[154] ^ m[155] ^ m[158] ^ m[159] ^ m[162] ^ m[163] ^ m[166] ^ m[167] ^ m[170] ^ m[171] ^ m[174] ^ m[176] ^ m[178] ^ m[180] ^ m[182] ^ m[185] ^ m[188] ^ m[191] ^ m[194] ^ m[195] ^ m[198] ^ m[201] ^ m[203] ^ m[205] ^ m[208] ^ m[209] ^ m[212] ^ m[215] ^ m[218] ^ m[221] ^ m[224] ^ m[225] ^ m[228] ^ m[231] ^ m[233] ^ m[235] ^ m[239] ^ m[241] ^ m[244] ^ m[245] ^ m[247] ^ m[252] ^ m[255] ^ m[258] ^ m[260] ^ m[262] ^ m[265] ^ m[268] ^ m[271] ^ m[274] ^ m[277] ^ m[279] ^ m[281] ^ m[284] ^ m[287] ^ m[289] ^ m[291] ^ m[293] ^ m[295] ^ m[297] ^ m[300] ^ m[302] ^ m[305] ^ m[307] ^ m[309] ^ m[311] ^ m[312] ^ m[315] ^ m[316] ^ m[319] ^ m[320] ^ m[323] ^ m[324] ^ m[327] ^ m[328] ^ m[331] ^ m[332] ^ m[335] ^ m[336] ^ m[339] ^ m[340] ^ m[343] ^ m[344] ^ m[347] ^ m[348] ^ m[351] ^ m[352] ^ m[355] ^ m[356] ^ m[359] ^ m[360] ^ m[363] ^ m[364] ^ m[367] ^ m[368] ^ m[371] ^ m[372] ^ m[375] ^ m[376] ^ m[379] ^ m[380] ^ m[383] ^ m[384] ^ m[387] ^ m[388] ^ m[390] ^ m[392] ^ m[394] ^ m[397] ^ m[398] ^ m[401] ^ m[402] ^ m[405] ^ m[406] ^ m[409] ^ m[410] ^ m[413] ^ m[414] ^ m[417] ^ m[418] ^ m[421] ^ m[422] ^ m[425] ^ m[426] ^ m[429] ^ m[430] ^ m[433] ^ m[434] ^ m[437] ^ m[438] ^ m[441] ^ m[442] ^ m[445] ^ m[446] ^ m[449] ^ m[450] ^ m[453] ^ m[454] ^ m[457] ^ m[459] ^ m[461] ^ m[463] ^ m[465] ^ m[467] ^ m[469] ^ m[471] ^ m[473] ^ m[475] ^ m[477] ^ m[479] ^ m[481] ^ m[483] ^ m[485] ^ m[487] ^ m[489] ^ m[491] ^ m[493] ^ m[495] ^ m[497] ^ m[499] ^ m[501] ^ m[503] ^ m[505] ^ m[507] ^ m[509] ^ m[511] ^ m[513] ^ m[515] ^ m[517] ^ m[519] ^ m[521] ^ m[523] ^ m[525] ^ m[527] ^ m[529] ^ m[531] ^ m[533] ^ m[535] ^ m[536] ^ m[539] ^ m[540] ^ m[543] ^ m[544] ^ m[547] ^ m[548] ^ m[551] ^ m[552] ^ m[555] ^ m[556] ^ m[557] ^ m[559] ^ m[561] ^ m[563] ^ m[565] ^ m[567] ^ m[569] ^ m[571] ^ m[573] ^ m[575] ^ m[577] ^ m[579] ^ m[581] ^ m[583] ^ m[585] ^ m[587] ^ m[589] ^ m[591] ^ m[593] ^ m[595] ^ m[597] ^ m[599] ^ m[601] ^ m[603] ^ m[605] ^ m[607] ^ m[609] ^ m[611] ^ m[613] ^ m[615] ^ m[617] ^ m[619] ^ m[621] ^ m[623] ^ m[625] ^ m[627] ^ m[629] ^ m[631] ^ m[633] ^ m[635] ^ m[637] ^ m[640] ^ m[641] ^ m[644] ^ m[645] ^ m[648] ^ m[649] ^ m[652] ^ m[653] ^ m[656] ^ m[657] ^ m[660] ^ m[661] ^ m[664] ^ m[665] ^ m[668] ^ m[669] ^ m[672] ^ m[673] ^ m[676] ^ m[677] ^ m[680] ^ m[681] ^ m[684] ^ m[685] ^ m[688] ^ m[689] ^ m[692] ^ m[693] ^ m[696] ^ m[697] ^ m[700] ^ m[701] ^ m[704] ^ m[705] ^ m[708] ^ m[710] ^ m[712] ^ m[714] ^ m[716] ^ m[718] ^ m[720] ^ m[722] ^ m[724] ^ m[726] ^ m[728] ^ m[730] ^ m[732] ^ m[734] ^ m[736] ^ m[738] ^ m[740] ^ m[742] ^ m[744] ^ m[746] ^ m[748] ^ m[750] ^ m[752] ^ m[754] ^ m[756] ^ m[758] ^ m[760] ^ m[762] ^ m[764] ^ m[766] ^ m[768] ^ m[770] ^ m[772] ^ m[774] ^ m[776] ^ m[778] ^ m[779] ^ m[782] ^ m[783] ^ m[786] ^ m[787] ^ m[790] ^ m[791] ^ m[794] ^ m[795] ^ m[798] ^ m[799] ^ m[802] ^ m[803] ^ m[806] ^ m[807] ^ m[810] ^ m[811] ^ m[813] ^ m[814] ^ m[816] ^ m[819] ^ m[820] ^ m[823] ^ m[824] ^ m[826] ^ m[827] ^ m[830] ^ m[831] ^ m[832] ^ m[834] ^ m[836] ^ m[838] ^ m[840] ^ m[841] ^ m[843] ^ m[844] ^ m[846] ^ m[848] ^ m[850] ^ m[852] ^ m[854] ^ m[856] ^ m[857] ^ m[859] ^ m[861] ^ m[862] ^ m[865] ^ m[866] ^ m[868] ^ m[869] ^ m[871] ^ m[872] ^ m[874] ^ m[876] ^ m[877] ^ m[878] ^ m[881] ^ m[883] ^ m[885] ^ m[886] ^ m[888] ^ m[891] ^ m[892] ^ m[893] ^ m[895] ^ m[898] ^ m[899] ^ m[901] ^ m[904] ^ m[905] ^ m[907] ^ m[909] ^ m[910] ^ m[913] ^ m[914] ^ m[916] ^ m[918] ^ m[920] ^ m[921] ^ m[922] ^ m[924] ^ m[926] ^ m[927] ^ m[930] ^ m[932] ^ m[934] ^ m[936] ^ m[937] ^ m[939] ^ m[941] ^ m[943] ^ m[945] ^ m[946] ^ m[948] ^ m[949] ^ m[951] ^ m[953] ^ m[954] ^ m[956] ^ m[959] ^ m[961] ^ m[962] ^ m[963] ^ m[964] ^ m[965] ^ m[966] ^ m[968] ^ m[971] ^ m[973] ^ m[974] ^ m[976] ^ m[977] ^ m[979] ^ m[982] ^ m[983] ^ m[985] ^ m[986] ^ m[989] ^ m[990] ^ m[992] ^ m[993] ^ m[995] ^ m[996] ^ m[997] ^ m[999] ^ m[1000] ^ m[1002] ^ m[1003] ^ m[1004] ^ m[1005] ^ m[1006] ^ m[1008] ^ m[1010] ^ m[1012];
    assign parity[8] = m[0] ^ m[1] ^ m[3] ^ m[6] ^ m[7] ^ m[10] ^ m[11] ^ m[14] ^ m[15] ^ m[18] ^ m[19] ^ m[22] ^ m[23] ^ m[26] ^ m[27] ^ m[30] ^ m[31] ^ m[34] ^ m[36] ^ m[37] ^ m[40] ^ m[41] ^ m[44] ^ m[45] ^ m[48] ^ m[49] ^ m[52] ^ m[53] ^ m[56] ^ m[57] ^ m[60] ^ m[61] ^ m[64] ^ m[65] ^ m[68] ^ m[70] ^ m[72] ^ m[74] ^ m[76] ^ m[78] ^ m[80] ^ m[82] ^ m[84] ^ m[86] ^ m[88] ^ m[90] ^ m[92] ^ m[94] ^ m[96] ^ m[98] ^ m[100] ^ m[102] ^ m[104] ^ m[106] ^ m[108] ^ m[110] ^ m[112] ^ m[114] ^ m[116] ^ m[118] ^ m[120] ^ m[122] ^ m[124] ^ m[126] ^ m[128] ^ m[130] ^ m[132] ^ m[134] ^ m[136] ^ m[138] ^ m[140] ^ m[142] ^ m[144] ^ m[146] ^ m[147] ^ m[150] ^ m[151] ^ m[154] ^ m[155] ^ m[158] ^ m[159] ^ m[162] ^ m[163] ^ m[166] ^ m[167] ^ m[170] ^ m[171] ^ m[174] ^ m[175] ^ m[178] ^ m[179] ^ m[181] ^ m[184] ^ m[187] ^ m[190] ^ m[193] ^ m[195] ^ m[197] ^ m[200] ^ m[202] ^ m[204] ^ m[207] ^ m[209] ^ m[211] ^ m[214] ^ m[217] ^ m[220] ^ m[223] ^ m[225] ^ m[227] ^ m[230] ^ m[232] ^ m[234] ^ m[237] ^ m[240] ^ m[243] ^ m[245] ^ m[248] ^ m[250] ^ m[253] ^ m[256] ^ m[258] ^ m[262] ^ m[265] ^ m[268] ^ m[271] ^ m[274] ^ m[277] ^ m[279] ^ m[281] ^ m[284] ^ m[287] ^ m[289] ^ m[291] ^ m[293] ^ m[295] ^ m[297] ^ m[300] ^ m[302] ^ m[304] ^ m[307] ^ m[309] ^ m[310] ^ m[312] ^ m[314] ^ m[316] ^ m[318] ^ m[320] ^ m[322] ^ m[324] ^ m[326] ^ m[328] ^ m[330] ^ m[332] ^ m[334] ^ m[336] ^ m[338] ^ m[340] ^ m[342] ^ m[344] ^ m[346] ^ m[348] ^ m[350] ^ m[352] ^ m[354] ^ m[356] ^ m[358] ^ m[360] ^ m[362] ^ m[364] ^ m[366] ^ m[368] ^ m[370] ^ m[372] ^ m[374] ^ m[376] ^ m[378] ^ m[380] ^ m[382] ^ m[384] ^ m[386] ^ m[388] ^ m[391] ^ m[392] ^ m[395] ^ m[396] ^ m[399] ^ m[400] ^ m[403] ^ m[404] ^ m[407] ^ m[408] ^ m[411] ^ m[412] ^ m[415] ^ m[416] ^ m[419] ^ m[420] ^ m[423] ^ m[424] ^ m[427] ^ m[428] ^ m[431] ^ m[432] ^ m[435] ^ m[436] ^ m[439] ^ m[440] ^ m[443] ^ m[444] ^ m[447] ^ m[448] ^ m[451] ^ m[452] ^ m[455] ^ m[456] ^ m[459] ^ m[460] ^ m[463] ^ m[464] ^ m[467] ^ m[468] ^ m[471] ^ m[472] ^ m[475] ^ m[476] ^ m[479] ^ m[480] ^ m[483] ^ m[484] ^ m[487] ^ m[488] ^ m[491] ^ m[492] ^ m[495] ^ m[496] ^ m[499] ^ m[500] ^ m[503] ^ m[504] ^ m[507] ^ m[508] ^ m[511] ^ m[512] ^ m[515] ^ m[516] ^ m[519] ^ m[520] ^ m[523] ^ m[524] ^ m[527] ^ m[528] ^ m[531] ^ m[532] ^ m[535] ^ m[537] ^ m[539] ^ m[541] ^ m[543] ^ m[545] ^ m[547] ^ m[549] ^ m[551] ^ m[553] ^ m[555] ^ m[556] ^ m[558] ^ m[559] ^ m[562] ^ m[563] ^ m[566] ^ m[567] ^ m[568] ^ m[571] ^ m[574] ^ m[575] ^ m[576] ^ m[579] ^ m[582] ^ m[583] ^ m[586] ^ m[587] ^ m[590] ^ m[591] ^ m[594] ^ m[595] ^ m[598] ^ m[599] ^ m[602] ^ m[603] ^ m[606] ^ m[607] ^ m[608] ^ m[611] ^ m[612] ^ m[615] ^ m[618] ^ m[619] ^ m[622] ^ m[623] ^ m[624] ^ m[627] ^ m[630] ^ m[631] ^ m[634] ^ m[635] ^ m[638] ^ m[639] ^ m[642] ^ m[643] ^ m[646] ^ m[647] ^ m[650] ^ m[651] ^ m[654] ^ m[655] ^ m[656] ^ m[659] ^ m[662] ^ m[663] ^ m[666] ^ m[667] ^ m[670] ^ m[671] ^ m[674] ^ m[675] ^ m[678] ^ m[679] ^ m[682] ^ m[683] ^ m[686] ^ m[687] ^ m[690] ^ m[691] ^ m[694] ^ m[695] ^ m[698] ^ m[699] ^ m[700] ^ m[703] ^ m[706] ^ m[707] ^ m[710] ^ m[711] ^ m[714] ^ m[715] ^ m[718] ^ m[719] ^ m[722] ^ m[723] ^ m[726] ^ m[727] ^ m[730] ^ m[731] ^ m[734] ^ m[735] ^ m[738] ^ m[739] ^ m[742] ^ m[743] ^ m[746] ^ m[747] ^ m[750] ^ m[751] ^ m[754] ^ m[755] ^ m[758] ^ m[759] ^ m[762] ^ m[763] ^ m[766] ^ m[767] ^ m[770] ^ m[771] ^ m[774] ^ m[775] ^ m[778] ^ m[780] ^ m[782] ^ m[784] ^ m[786] ^ m[788] ^ m[790] ^ m[792] ^ m[794] ^ m[796] ^ m[798] ^ m[800] ^ m[802] ^ m[804] ^ m[806] ^ m[808] ^ m[810] ^ m[812] ^ m[814] ^ m[816] ^ m[818] ^ m[819] ^ m[821] ^ m[823] ^ m[825] ^ m[826] ^ m[827] ^ m[829] ^ m[832] ^ m[833] ^ m[835] ^ m[837] ^ m[839] ^ m[840] ^ m[841] ^ m[843] ^ m[845] ^ m[847] ^ m[850] ^ m[851] ^ m[853] ^ m[855] ^ m[857] ^ m[859] ^ m[860] ^ m[862] ^ m[864] ^ m[865] ^ m[867] ^ m[868] ^ m[869] ^ m[871] ^ m[873] ^ m[874] ^ m[875] ^ m[878] ^ m[880] ^ m[883] ^ m[884] ^ m[886] ^ m[888] ^ m[889] ^ m[891] ^ m[893] ^ m[895] ^ m[896] ^ m[898] ^ m[900] ^ m[901] ^ m[902] ^ m[904] ^ m[907] ^ m[909] ^ m[910] ^ m[911] ^ m[913] ^ m[916] ^ m[918] ^ m[920] ^ m[921] ^ m[922] ^ m[924] ^ m[926] ^ m[929] ^ m[930] ^ m[932] ^ m[934] ^ m[936] ^ m[937] ^ m[939] ^ m[941] ^ m[943] ^ m[945] ^ m[946] ^ m[948] ^ m[949] ^ m[951] ^ m[953] ^ m[954] ^ m[957] ^ m[959] ^ m[961] ^ m[962] ^ m[963] ^ m[965] ^ m[966] ^ m[968] ^ m[969] ^ m[971] ^ m[972] ^ m[974] ^ m[975] ^ m[976] ^ m[977] ^ m[979] ^ m[980] ^ m[981] ^ m[982] ^ m[984] ^ m[985] ^ m[987] ^ m[988] ^ m[989] ^ m[991] ^ m[992] ^ m[994] ^ m[996] ^ m[997] ^ m[999] ^ m[1003] ^ m[1004] ^ m[1006] ^ m[1007] ^ m[1009] ^ m[1012];
    assign parity[9] = m[0] ^ m[1] ^ m[3] ^ m[5] ^ m[7] ^ m[9] ^ m[11] ^ m[13] ^ m[15] ^ m[17] ^ m[19] ^ m[21] ^ m[23] ^ m[25] ^ m[27] ^ m[29] ^ m[31] ^ m[33] ^ m[35] ^ m[38] ^ m[39] ^ m[42] ^ m[43] ^ m[46] ^ m[47] ^ m[50] ^ m[51] ^ m[54] ^ m[55] ^ m[58] ^ m[59] ^ m[62] ^ m[63] ^ m[66] ^ m[67] ^ m[70] ^ m[71] ^ m[74] ^ m[75] ^ m[78] ^ m[79] ^ m[82] ^ m[83] ^ m[86] ^ m[87] ^ m[90] ^ m[91] ^ m[94] ^ m[95] ^ m[98] ^ m[99] ^ m[102] ^ m[103] ^ m[106] ^ m[107] ^ m[110] ^ m[111] ^ m[114] ^ m[115] ^ m[118] ^ m[119] ^ m[122] ^ m[123] ^ m[126] ^ m[127] ^ m[130] ^ m[131] ^ m[134] ^ m[135] ^ m[138] ^ m[139] ^ m[142] ^ m[143] ^ m[146] ^ m[148] ^ m[150] ^ m[152] ^ m[154] ^ m[156] ^ m[158] ^ m[160] ^ m[162] ^ m[164] ^ m[166] ^ m[168] ^ m[170] ^ m[172] ^ m[174] ^ m[176] ^ m[178] ^ m[180] ^ m[183] ^ m[186] ^ m[189] ^ m[192] ^ m[195] ^ m[197] ^ m[199] ^ m[202] ^ m[204] ^ m[206] ^ m[209] ^ m[211] ^ m[213] ^ m[216] ^ m[219] ^ m[222] ^ m[225] ^ m[227] ^ m[229] ^ m[232] ^ m[234] ^ m[236] ^ m[239] ^ m[242] ^ m[245] ^ m[247] ^ m[249] ^ m[252] ^ m[255] ^ m[258] ^ m[260] ^ m[262] ^ m[265] ^ m[268] ^ m[271] ^ m[274] ^ m[277] ^ m[279] ^ m[281] ^ m[284] ^ m[287] ^ m[289] ^ m[291] ^ m[293] ^ m[294] ^ m[297] ^ m[298] ^ m[302] ^ m[304] ^ m[305] ^ m[309] ^ m[310] ^ m[312] ^ m[314] ^ m[316] ^ m[318] ^ m[320] ^ m[322] ^ m[324] ^ m[326] ^ m[328] ^ m[330] ^ m[332] ^ m[334] ^ m[336] ^ m[338] ^ m[340] ^ m[342] ^ m[344] ^ m[346] ^ m[348] ^ m[350] ^ m[352] ^ m[354] ^ m[356] ^ m[358] ^ m[360] ^ m[362] ^ m[364] ^ m[366] ^ m[368] ^ m[370] ^ m[372] ^ m[374] ^ m[376] ^ m[378] ^ m[380] ^ m[382] ^ m[384] ^ m[386] ^ m[388] ^ m[390] ^ m[392] ^ m[394] ^ m[396] ^ m[398] ^ m[400] ^ m[402] ^ m[404] ^ m[406] ^ m[408] ^ m[410] ^ m[412] ^ m[414] ^ m[416] ^ m[418] ^ m[420] ^ m[422] ^ m[424] ^ m[426] ^ m[428] ^ m[430] ^ m[432] ^ m[434] ^ m[436] ^ m[438] ^ m[440] ^ m[442] ^ m[444] ^ m[446] ^ m[448] ^ m[450] ^ m[452] ^ m[454] ^ m[456] ^ m[458] ^ m[460] ^ m[462] ^ m[464] ^ m[466] ^ m[468] ^ m[470] ^ m[472] ^ m[474] ^ m[476] ^ m[478] ^ m[480] ^ m[482] ^ m[484] ^ m[486] ^ m[488] ^ m[490] ^ m[492] ^ m[494] ^ m[496] ^ m[498] ^ m[500] ^ m[502] ^ m[504] ^ m[506] ^ m[508] ^ m[510] ^ m[512] ^ m[514] ^ m[516] ^ m[518] ^ m[520] ^ m[522] ^ m[524] ^ m[526] ^ m[528] ^ m[530] ^ m[532] ^ m[534] ^ m[536] ^ m[538] ^ m[540] ^ m[542] ^ m[544] ^ m[546] ^ m[548] ^ m[550] ^ m[552] ^ m[554] ^ m[555] ^ m[558] ^ m[560] ^ m[561] ^ m[564] ^ m[565] ^ m[568] ^ m[570] ^ m[572] ^ m[573] ^ m[576] ^ m[578] ^ m[580] ^ m[581] ^ m[584] ^ m[585] ^ m[588] ^ m[589] ^ m[592] ^ m[593] ^ m[596] ^ m[597] ^ m[600] ^ m[601] ^ m[604] ^ m[605] ^ m[608] ^ m[610] ^ m[612] ^ m[614] ^ m[616] ^ m[617] ^ m[620] ^ m[621] ^ m[624] ^ m[626] ^ m[628] ^ m[629] ^ m[632] ^ m[633] ^ m[636] ^ m[637] ^ m[640] ^ m[641] ^ m[644] ^ m[645] ^ m[648] ^ m[649] ^ m[652] ^ m[653] ^ m[656] ^ m[658] ^ m[660] ^ m[661] ^ m[664] ^ m[665] ^ m[668] ^ m[669] ^ m[672] ^ m[673] ^ m[676] ^ m[677] ^ m[680] ^ m[681] ^ m[684] ^ m[685] ^ m[688] ^ m[689] ^ m[692] ^ m[693] ^ m[696] ^ m[697] ^ m[700] ^ m[702] ^ m[704] ^ m[705] ^ m[708] ^ m[709] ^ m[712] ^ m[713] ^ m[716] ^ m[717] ^ m[720] ^ m[721] ^ m[724] ^ m[725] ^ m[728] ^ m[729] ^ m[732] ^ m[733] ^ m[736] ^ m[737] ^ m[740] ^ m[741] ^ m[744] ^ m[745] ^ m[748] ^ m[749] ^ m[752] ^ m[753] ^ m[756] ^ m[757] ^ m[760] ^ m[761] ^ m[764] ^ m[765] ^ m[768] ^ m[769] ^ m[772] ^ m[773] ^ m[776] ^ m[777] ^ m[780] ^ m[781] ^ m[784] ^ m[785] ^ m[788] ^ m[789] ^ m[792] ^ m[793] ^ m[796] ^ m[797] ^ m[800] ^ m[801] ^ m[804] ^ m[805] ^ m[808] ^ m[809] ^ m[812] ^ m[814] ^ m[815] ^ m[818] ^ m[819] ^ m[821] ^ m[822] ^ m[825] ^ m[827] ^ m[829] ^ m[830] ^ m[832] ^ m[833] ^ m[835] ^ m[837] ^ m[839] ^ m[841] ^ m[843] ^ m[845] ^ m[847] ^ m[848] ^ m[850] ^ m[851] ^ m[853] ^ m[855] ^ m[857] ^ m[859] ^ m[860] ^ m[862] ^ m[864] ^ m[865] ^ m[867] ^ m[869] ^ m[871] ^ m[873] ^ m[875] ^ m[876] ^ m[878] ^ m[880] ^ m[881] ^ m[883] ^ m[884] ^ m[886] ^ m[888] ^ m[889] ^ m[891] ^ m[893] ^ m[895] ^ m[896] ^ m[898] ^ m[900] ^ m[902] ^ m[904] ^ m[905] ^ m[907] ^ m[909] ^ m[911] ^ m[913] ^ m[914] ^ m[916] ^ m[918] ^ m[920] ^ m[922] ^ m[924] ^ m[926] ^ m[927] ^ m[929] ^ m[930] ^ m[932] ^ m[934] ^ m[936] ^ m[937] ^ m[939] ^ m[941] ^ m[943] ^ m[945] ^ m[946] ^ m[948] ^ m[949] ^ m[951] ^ m[953] ^ m[954] ^ m[956] ^ m[957] ^ m[959] ^ m[962] ^ m[963] ^ m[964] ^ m[965] ^ m[966] ^ m[968] ^ m[969] ^ m[971] ^ m[973] ^ m[974] ^ m[976] ^ m[977] ^ m[979] ^ m[980] ^ m[981] ^ m[983] ^ m[984] ^ m[986] ^ m[987] ^ m[988] ^ m[990] ^ m[991] ^ m[993] ^ m[994] ^ m[995] ^ m[999] ^ m[1000] ^ m[1002] ^ m[1004] ^ m[1005] ^ m[1008] ^ m[1010] ^ m[1012];
    assign parity[10] = m[0] ^ m[1] ^ m[2] ^ m[5] ^ m[6] ^ m[9] ^ m[10] ^ m[13] ^ m[14] ^ m[17] ^ m[18] ^ m[21] ^ m[22] ^ m[25] ^ m[26] ^ m[29] ^ m[30] ^ m[33] ^ m[34] ^ m[37] ^ m[38] ^ m[41] ^ m[42] ^ m[45] ^ m[46] ^ m[49] ^ m[50] ^ m[53] ^ m[54] ^ m[57] ^ m[58] ^ m[61] ^ m[62] ^ m[65] ^ m[66] ^ m[69] ^ m[70] ^ m[73] ^ m[74] ^ m[77] ^ m[78] ^ m[81] ^ m[82] ^ m[85] ^ m[86] ^ m[89] ^ m[90] ^ m[93] ^ m[94] ^ m[97] ^ m[98] ^ m[101] ^ m[102] ^ m[105] ^ m[106] ^ m[109] ^ m[110] ^ m[113] ^ m[114] ^ m[117] ^ m[118] ^ m[121] ^ m[122] ^ m[125] ^ m[126] ^ m[129] ^ m[130] ^ m[133] ^ m[134] ^ m[137] ^ m[138] ^ m[141] ^ m[142] ^ m[145] ^ m[146] ^ m[149] ^ m[150] ^ m[153] ^ m[154] ^ m[157] ^ m[158] ^ m[161] ^ m[162] ^ m[165] ^ m[166] ^ m[169] ^ m[170] ^ m[173] ^ m[174] ^ m[177] ^ m[178] ^ m[183] ^ m[186] ^ m[189] ^ m[192] ^ m[195] ^ m[197] ^ m[199] ^ m[202] ^ m[204] ^ m[206] ^ m[209] ^ m[211] ^ m[213] ^ m[216] ^ m[219] ^ m[222] ^ m[225] ^ m[227] ^ m[229] ^ m[232] ^ m[234] ^ m[236] ^ m[239] ^ m[242] ^ m[245] ^ m[247] ^ m[249] ^ m[252] ^ m[255] ^ m[258] ^ m[260] ^ m[262] ^ m[265] ^ m[268] ^ m[271] ^ m[274] ^ m[277] ^ m[279] ^ m[281] ^ m[284] ^ m[287] ^ m[289] ^ m[291] ^ m[293] ^ m[294] ^ m[297] ^ m[298] ^ m[300] ^ m[304] ^ m[305] ^ m[307] ^ m[310] ^ m[311] ^ m[314] ^ m[315] ^ m[318] ^ m[319] ^ m[322] ^ m[323] ^ m[326] ^ m[327] ^ m[330] ^ m[331] ^ m[334] ^ m[335] ^ m[338] ^ m[339] ^ m[342] ^ m[343] ^ m[346] ^ m[347] ^ m[350] ^ m[351] ^ m[354] ^ m[355] ^ m[358] ^ m[359] ^ m[362] ^ m[363] ^ m[366] ^ m[367] ^ m[370] ^ m[371] ^ m[374] ^ m[375] ^ m[378] ^ m[379] ^ m[382] ^ m[383] ^ m[386] ^ m[387] ^ m[390] ^ m[391] ^ m[394] ^ m[395] ^ m[398] ^ m[399] ^ m[402] ^ m[403] ^ m[406] ^ m[407] ^ m[410] ^ m[411] ^ m[414] ^ m[415] ^ m[418] ^ m[419] ^ m[422] ^ m[423] ^ m[426] ^ m[427] ^ m[430] ^ m[431] ^ m[434] ^ m[435] ^ m[438] ^ m[439] ^ m[442] ^ m[443] ^ m[446] ^ m[447] ^ m[450] ^ m[451] ^ m[454] ^ m[455] ^ m[458] ^ m[459] ^ m[462] ^ m[463] ^ m[466] ^ m[467] ^ m[470] ^ m[471] ^ m[474] ^ m[475] ^ m[478] ^ m[479] ^ m[482] ^ m[483] ^ m[486] ^ m[487] ^ m[490] ^ m[491] ^ m[494] ^ m[495] ^ m[498] ^ m[499] ^ m[502] ^ m[503] ^ m[506] ^ m[507] ^ m[510] ^ m[511] ^ m[514] ^ m[515] ^ m[518] ^ m[519] ^ m[522] ^ m[523] ^ m[526] ^ m[527] ^ m[530] ^ m[531] ^ m[534] ^ m[535] ^ m[538] ^ m[539] ^ m[542] ^ m[543] ^ m[546] ^ m[547] ^ m[550] ^ m[551] ^ m[554] ^ m[556] ^ m[557] ^ m[559] ^ m[560] ^ m[563] ^ m[564] ^ m[567] ^ m[569] ^ m[571] ^ m[572] ^ m[575] ^ m[577] ^ m[579] ^ m[580] ^ m[583] ^ m[584] ^ m[587] ^ m[588] ^ m[591] ^ m[592] ^ m[595] ^ m[596] ^ m[599] ^ m[600] ^ m[603] ^ m[604] ^ m[607] ^ m[609] ^ m[611] ^ m[613] ^ m[615] ^ m[616] ^ m[619] ^ m[620] ^ m[623] ^ m[625] ^ m[627] ^ m[628] ^ m[631] ^ m[632] ^ m[635] ^ m[636] ^ m[639] ^ m[640] ^ m[643] ^ m[644] ^ m[647] ^ m[648] ^ m[651] ^ m[652] ^ m[655] ^ m[657] ^ m[659] ^ m[660] ^ m[663] ^ m[664] ^ m[667] ^ m[668] ^ m[671] ^ m[672] ^ m[675] ^ m[676] ^ m[679] ^ m[680] ^ m[683] ^ m[684] ^ m[687] ^ m[688] ^ m[691] ^ m[692] ^ m[695] ^ m[696] ^ m[699] ^ m[701] ^ m[703] ^ m[704] ^ m[707] ^ m[708] ^ m[711] ^ m[712] ^ m[715] ^ m[716] ^ m[719] ^ m[720] ^ m[723] ^ m[724] ^ m[727] ^ m[728] ^ m[731] ^ m[732] ^ m[735] ^ m[736] ^ m[739] ^ m[740] ^ m[743] ^ m[744] ^ m[747] ^ m[748] ^ m[751] ^ m[752] ^ m[755] ^ m[756] ^ m[759] ^ m[760] ^ m[763] ^ m[764] ^ m[767] ^ m[768] ^ m[771] ^ m[772] ^ m[775] ^ m[776] ^ m[779] ^ m[780] ^ m[783] ^ m[784] ^ m[787] ^ m[788] ^ m[791] ^ m[792] ^ m[795] ^ m[796] ^ m[799] ^ m[800] ^ m[803] ^ m[804] ^ m[807] ^ m[808] ^ m[811] ^ m[813] ^ m[814] ^ m[817] ^ m[818] ^ m[820] ^ m[821] ^ m[824] ^ m[825] ^ m[828] ^ m[829] ^ m[831] ^ m[832] ^ m[834] ^ m[836] ^ m[838] ^ m[839] ^ m[842] ^ m[843] ^ m[844] ^ m[846] ^ m[849] ^ m[850] ^ m[852] ^ m[854] ^ m[856] ^ m[858] ^ m[859] ^ m[861] ^ m[863] ^ m[864] ^ m[866] ^ m[867] ^ m[870] ^ m[871] ^ m[872] ^ m[873] ^ m[875] ^ m[877] ^ m[879] ^ m[882] ^ m[883] ^ m[885] ^ m[887] ^ m[888] ^ m[890] ^ m[892] ^ m[894] ^ m[895] ^ m[897] ^ m[899] ^ m[900] ^ m[903] ^ m[904] ^ m[906] ^ m[908] ^ m[909] ^ m[912] ^ m[913] ^ m[915] ^ m[917] ^ m[919] ^ m[920] ^ m[922] ^ m[923] ^ m[925] ^ m[928] ^ m[929] ^ m[931] ^ m[933] ^ m[935] ^ m[936] ^ m[938] ^ m[940] ^ m[942] ^ m[944] ^ m[945] ^ m[947] ^ m[949] ^ m[950] ^ m[952] ^ m[954] ^ m[955] ^ m[957] ^ m[958] ^ m[960] ^ m[961] ^ m[963] ^ m[965] ^ m[966] ^ m[967] ^ m[969] ^ m[970] ^ m[972] ^ m[974] ^ m[975] ^ m[977] ^ m[978] ^ m[980] ^ m[981] ^ m[982] ^ m[984] ^ m[985] ^ m[987] ^ m[988] ^ m[989] ^ m[991] ^ m[992] ^ m[994] ^ m[996] ^ m[997] ^ m[998] ^ m[1001] ^ m[1003] ^ m[1006] ^ m[1007] ^ m[1009] ^ m[1011];
  end else if ((CodewordWidth == 2048) && (MessageWidth == 2036)) begin : gen_2048_2036
    `BR_ASSERT_STATIC(parity_width_matches_a, ParityWidth == 12)
    assign parity[0] = m[1] ^ m[3] ^ m[5] ^ m[7] ^ m[9] ^ m[11] ^ m[13] ^ m[15] ^ m[17] ^ m[18] ^ m[21] ^ m[23] ^ m[25] ^ m[27] ^ m[29] ^ m[31] ^ m[33] ^ m[35] ^ m[36] ^ m[39] ^ m[41] ^ m[43] ^ m[45] ^ m[47] ^ m[49] ^ m[51] ^ m[52] ^ m[55] ^ m[57] ^ m[59] ^ m[61] ^ m[63] ^ m[65] ^ m[66] ^ m[69] ^ m[71] ^ m[73] ^ m[75] ^ m[77] ^ m[78] ^ m[81] ^ m[83] ^ m[85] ^ m[87] ^ m[88] ^ m[91] ^ m[93] ^ m[95] ^ m[96] ^ m[99] ^ m[101] ^ m[102] ^ m[105] ^ m[106] ^ m[108] ^ m[111] ^ m[113] ^ m[115] ^ m[117] ^ m[119] ^ m[121] ^ m[123] ^ m[125] ^ m[126] ^ m[129] ^ m[131] ^ m[133] ^ m[135] ^ m[137] ^ m[139] ^ m[141] ^ m[142] ^ m[145] ^ m[147] ^ m[149] ^ m[151] ^ m[153] ^ m[155] ^ m[156] ^ m[159] ^ m[161] ^ m[163] ^ m[165] ^ m[167] ^ m[168] ^ m[171] ^ m[173] ^ m[175] ^ m[177] ^ m[178] ^ m[181] ^ m[183] ^ m[185] ^ m[186] ^ m[189] ^ m[191] ^ m[192] ^ m[195] ^ m[196] ^ m[198] ^ m[201] ^ m[203] ^ m[205] ^ m[207] ^ m[209] ^ m[211] ^ m[213] ^ m[214] ^ m[217] ^ m[219] ^ m[221] ^ m[223] ^ m[225] ^ m[227] ^ m[228] ^ m[231] ^ m[233] ^ m[235] ^ m[237] ^ m[239] ^ m[240] ^ m[243] ^ m[245] ^ m[247] ^ m[249] ^ m[250] ^ m[253] ^ m[255] ^ m[257] ^ m[258] ^ m[261] ^ m[263] ^ m[264] ^ m[267] ^ m[268] ^ m[270] ^ m[273] ^ m[275] ^ m[277] ^ m[279] ^ m[281] ^ m[283] ^ m[284] ^ m[287] ^ m[289] ^ m[291] ^ m[293] ^ m[295] ^ m[296] ^ m[299] ^ m[301] ^ m[303] ^ m[305] ^ m[306] ^ m[309] ^ m[311] ^ m[313] ^ m[314] ^ m[317] ^ m[319] ^ m[320] ^ m[323] ^ m[324] ^ m[326] ^ m[329] ^ m[331] ^ m[333] ^ m[335] ^ m[337] ^ m[338] ^ m[341] ^ m[343] ^ m[345] ^ m[347] ^ m[348] ^ m[351] ^ m[353] ^ m[355] ^ m[356] ^ m[359] ^ m[361] ^ m[362] ^ m[365] ^ m[366] ^ m[368] ^ m[371] ^ m[373] ^ m[375] ^ m[377] ^ m[378] ^ m[381] ^ m[383] ^ m[385] ^ m[386] ^ m[389] ^ m[391] ^ m[392] ^ m[395] ^ m[396] ^ m[398] ^ m[401] ^ m[403] ^ m[405] ^ m[406] ^ m[409] ^ m[411] ^ m[412] ^ m[415] ^ m[416] ^ m[418] ^ m[421] ^ m[423] ^ m[424] ^ m[427] ^ m[428] ^ m[430] ^ m[433] ^ m[434] ^ m[436] ^ m[438] ^ m[441] ^ m[443] ^ m[445] ^ m[447] ^ m[449] ^ m[451] ^ m[453] ^ m[454] ^ m[457] ^ m[459] ^ m[461] ^ m[463] ^ m[465] ^ m[467] ^ m[468] ^ m[471] ^ m[473] ^ m[475] ^ m[477] ^ m[479] ^ m[480] ^ m[483] ^ m[485] ^ m[487] ^ m[489] ^ m[490] ^ m[493] ^ m[495] ^ m[497] ^ m[498] ^ m[501] ^ m[503] ^ m[504] ^ m[507] ^ m[508] ^ m[510] ^ m[513] ^ m[515] ^ m[517] ^ m[519] ^ m[521] ^ m[523] ^ m[524] ^ m[527] ^ m[529] ^ m[531] ^ m[533] ^ m[535] ^ m[536] ^ m[539] ^ m[541] ^ m[543] ^ m[545] ^ m[546] ^ m[549] ^ m[551] ^ m[553] ^ m[554] ^ m[557] ^ m[559] ^ m[560] ^ m[563] ^ m[564] ^ m[566] ^ m[569] ^ m[571] ^ m[573] ^ m[575] ^ m[577] ^ m[578] ^ m[581] ^ m[583] ^ m[585] ^ m[587] ^ m[588] ^ m[591] ^ m[593] ^ m[595] ^ m[596] ^ m[599] ^ m[601] ^ m[602] ^ m[605] ^ m[606] ^ m[608] ^ m[611] ^ m[613] ^ m[615] ^ m[617] ^ m[618] ^ m[621] ^ m[623] ^ m[625] ^ m[626] ^ m[629] ^ m[631] ^ m[632] ^ m[635] ^ m[636] ^ m[638] ^ m[641] ^ m[643] ^ m[645] ^ m[646] ^ m[649] ^ m[651] ^ m[652] ^ m[655] ^ m[656] ^ m[658] ^ m[661] ^ m[663] ^ m[664] ^ m[667] ^ m[668] ^ m[670] ^ m[673] ^ m[674] ^ m[676] ^ m[678] ^ m[681] ^ m[683] ^ m[685] ^ m[687] ^ m[689] ^ m[691] ^ m[692] ^ m[695] ^ m[697] ^ m[699] ^ m[701] ^ m[703] ^ m[704] ^ m[707] ^ m[709] ^ m[711] ^ m[713] ^ m[714] ^ m[717] ^ m[719] ^ m[721] ^ m[722] ^ m[725] ^ m[727] ^ m[728] ^ m[731] ^ m[732] ^ m[734] ^ m[737] ^ m[739] ^ m[741] ^ m[743] ^ m[745] ^ m[746] ^ m[749] ^ m[751] ^ m[753] ^ m[755] ^ m[756] ^ m[759] ^ m[761] ^ m[763] ^ m[764] ^ m[767] ^ m[769] ^ m[770] ^ m[773] ^ m[774] ^ m[776] ^ m[779] ^ m[781] ^ m[783] ^ m[785] ^ m[786] ^ m[789] ^ m[791] ^ m[793] ^ m[794] ^ m[797] ^ m[799] ^ m[800] ^ m[803] ^ m[804] ^ m[806] ^ m[809] ^ m[811] ^ m[813] ^ m[814] ^ m[817] ^ m[819] ^ m[820] ^ m[823] ^ m[824] ^ m[826] ^ m[829] ^ m[831] ^ m[832] ^ m[835] ^ m[836] ^ m[838] ^ m[841] ^ m[842] ^ m[844] ^ m[846] ^ m[849] ^ m[851] ^ m[853] ^ m[855] ^ m[857] ^ m[858] ^ m[861] ^ m[863] ^ m[865] ^ m[867] ^ m[868] ^ m[871] ^ m[873] ^ m[875] ^ m[876] ^ m[879] ^ m[881] ^ m[882] ^ m[885] ^ m[886] ^ m[888] ^ m[891] ^ m[893] ^ m[895] ^ m[897] ^ m[898] ^ m[901] ^ m[903] ^ m[905] ^ m[906] ^ m[909] ^ m[911] ^ m[912] ^ m[915] ^ m[916] ^ m[918] ^ m[921] ^ m[923] ^ m[925] ^ m[926] ^ m[929] ^ m[931] ^ m[932] ^ m[935] ^ m[936] ^ m[938] ^ m[941] ^ m[943] ^ m[944] ^ m[947] ^ m[948] ^ m[950] ^ m[953] ^ m[954] ^ m[956] ^ m[958] ^ m[961] ^ m[963] ^ m[965] ^ m[967] ^ m[968] ^ m[971] ^ m[973] ^ m[975] ^ m[976] ^ m[979] ^ m[981] ^ m[982] ^ m[985] ^ m[986] ^ m[988] ^ m[991] ^ m[993] ^ m[995] ^ m[996] ^ m[999] ^ m[1001] ^ m[1002] ^ m[1005] ^ m[1006] ^ m[1008] ^ m[1011] ^ m[1013] ^ m[1014] ^ m[1017] ^ m[1018] ^ m[1020] ^ m[1023] ^ m[1024] ^ m[1026] ^ m[1028] ^ m[1031] ^ m[1033] ^ m[1035] ^ m[1036] ^ m[1039] ^ m[1041] ^ m[1042] ^ m[1045] ^ m[1046] ^ m[1048] ^ m[1051] ^ m[1053] ^ m[1054] ^ m[1057] ^ m[1058] ^ m[1060] ^ m[1063] ^ m[1064] ^ m[1066] ^ m[1068] ^ m[1071] ^ m[1073] ^ m[1074] ^ m[1077] ^ m[1078] ^ m[1080] ^ m[1083] ^ m[1084] ^ m[1086] ^ m[1088] ^ m[1091] ^ m[1092] ^ m[1094] ^ m[1096] ^ m[1098] ^ m[1101] ^ m[1103] ^ m[1105] ^ m[1107] ^ m[1109] ^ m[1111] ^ m[1112] ^ m[1115] ^ m[1117] ^ m[1119] ^ m[1121] ^ m[1123] ^ m[1124] ^ m[1127] ^ m[1129] ^ m[1131] ^ m[1133] ^ m[1134] ^ m[1137] ^ m[1139] ^ m[1141] ^ m[1142] ^ m[1145] ^ m[1147] ^ m[1148] ^ m[1151] ^ m[1152] ^ m[1154] ^ m[1157] ^ m[1159] ^ m[1161] ^ m[1163] ^ m[1165] ^ m[1166] ^ m[1169] ^ m[1171] ^ m[1173] ^ m[1175] ^ m[1176] ^ m[1179] ^ m[1181] ^ m[1183] ^ m[1184] ^ m[1187] ^ m[1189] ^ m[1190] ^ m[1193] ^ m[1194] ^ m[1196] ^ m[1199] ^ m[1201] ^ m[1203] ^ m[1205] ^ m[1206] ^ m[1209] ^ m[1211] ^ m[1213] ^ m[1214] ^ m[1217] ^ m[1219] ^ m[1220] ^ m[1223] ^ m[1224] ^ m[1226] ^ m[1229] ^ m[1231] ^ m[1233] ^ m[1234] ^ m[1237] ^ m[1239] ^ m[1240] ^ m[1243] ^ m[1244] ^ m[1246] ^ m[1249] ^ m[1251] ^ m[1252] ^ m[1255] ^ m[1256] ^ m[1258] ^ m[1261] ^ m[1262] ^ m[1264] ^ m[1266] ^ m[1269] ^ m[1271] ^ m[1273] ^ m[1275] ^ m[1277] ^ m[1278] ^ m[1281] ^ m[1283] ^ m[1285] ^ m[1287] ^ m[1288] ^ m[1291] ^ m[1293] ^ m[1295] ^ m[1296] ^ m[1299] ^ m[1301] ^ m[1302] ^ m[1305] ^ m[1306] ^ m[1308] ^ m[1311] ^ m[1313] ^ m[1315] ^ m[1317] ^ m[1318] ^ m[1321] ^ m[1323] ^ m[1325] ^ m[1326] ^ m[1329] ^ m[1331] ^ m[1332] ^ m[1335] ^ m[1336] ^ m[1338] ^ m[1341] ^ m[1343] ^ m[1345] ^ m[1346] ^ m[1349] ^ m[1351] ^ m[1352] ^ m[1355] ^ m[1356] ^ m[1358] ^ m[1361] ^ m[1363] ^ m[1364] ^ m[1367] ^ m[1368] ^ m[1370] ^ m[1373] ^ m[1374] ^ m[1376] ^ m[1378] ^ m[1381] ^ m[1383] ^ m[1385] ^ m[1387] ^ m[1388] ^ m[1391] ^ m[1393] ^ m[1395] ^ m[1396] ^ m[1399] ^ m[1401] ^ m[1402] ^ m[1405] ^ m[1406] ^ m[1408] ^ m[1411] ^ m[1413] ^ m[1415] ^ m[1416] ^ m[1419] ^ m[1421] ^ m[1422] ^ m[1425] ^ m[1426] ^ m[1428] ^ m[1431] ^ m[1433] ^ m[1434] ^ m[1437] ^ m[1438] ^ m[1440] ^ m[1443] ^ m[1444] ^ m[1446] ^ m[1448] ^ m[1451] ^ m[1453] ^ m[1455] ^ m[1456] ^ m[1459] ^ m[1461] ^ m[1462] ^ m[1465] ^ m[1466] ^ m[1468] ^ m[1471] ^ m[1473] ^ m[1474] ^ m[1477] ^ m[1478] ^ m[1480] ^ m[1483] ^ m[1484] ^ m[1486] ^ m[1488] ^ m[1491] ^ m[1493] ^ m[1494] ^ m[1497] ^ m[1498] ^ m[1500] ^ m[1503] ^ m[1504] ^ m[1506] ^ m[1508] ^ m[1511] ^ m[1512] ^ m[1514] ^ m[1516] ^ m[1518] ^ m[1521] ^ m[1523] ^ m[1525] ^ m[1527] ^ m[1529] ^ m[1530] ^ m[1533] ^ m[1535] ^ m[1537] ^ m[1539] ^ m[1540] ^ m[1543] ^ m[1545] ^ m[1547] ^ m[1548] ^ m[1551] ^ m[1553] ^ m[1554] ^ m[1557] ^ m[1558] ^ m[1560] ^ m[1563] ^ m[1565] ^ m[1567] ^ m[1569] ^ m[1570] ^ m[1573] ^ m[1575] ^ m[1577] ^ m[1578] ^ m[1581] ^ m[1583] ^ m[1584] ^ m[1587] ^ m[1588] ^ m[1590] ^ m[1593] ^ m[1595] ^ m[1597] ^ m[1598] ^ m[1601] ^ m[1603] ^ m[1604] ^ m[1607] ^ m[1608] ^ m[1610] ^ m[1613] ^ m[1615] ^ m[1616] ^ m[1619] ^ m[1620] ^ m[1622] ^ m[1625] ^ m[1626] ^ m[1628] ^ m[1630] ^ m[1633] ^ m[1635] ^ m[1637] ^ m[1639] ^ m[1640] ^ m[1643] ^ m[1645] ^ m[1647] ^ m[1648] ^ m[1651] ^ m[1653] ^ m[1654] ^ m[1657] ^ m[1658] ^ m[1660] ^ m[1663] ^ m[1665] ^ m[1667] ^ m[1668] ^ m[1671] ^ m[1673] ^ m[1674] ^ m[1677] ^ m[1678] ^ m[1680] ^ m[1683] ^ m[1685] ^ m[1686] ^ m[1689] ^ m[1690] ^ m[1692] ^ m[1695] ^ m[1696] ^ m[1698] ^ m[1700] ^ m[1703] ^ m[1705] ^ m[1707] ^ m[1708] ^ m[1711] ^ m[1713] ^ m[1714] ^ m[1717] ^ m[1718] ^ m[1720] ^ m[1723] ^ m[1725] ^ m[1726] ^ m[1729] ^ m[1730] ^ m[1732] ^ m[1735] ^ m[1736] ^ m[1738] ^ m[1740] ^ m[1743] ^ m[1745] ^ m[1746] ^ m[1749] ^ m[1750] ^ m[1752] ^ m[1755] ^ m[1756] ^ m[1758] ^ m[1760] ^ m[1763] ^ m[1764] ^ m[1766] ^ m[1768] ^ m[1770] ^ m[1773] ^ m[1775] ^ m[1777] ^ m[1779] ^ m[1780] ^ m[1783] ^ m[1785] ^ m[1787] ^ m[1788] ^ m[1791] ^ m[1793] ^ m[1794] ^ m[1797] ^ m[1798] ^ m[1800] ^ m[1803] ^ m[1805] ^ m[1807] ^ m[1808] ^ m[1811] ^ m[1813] ^ m[1814] ^ m[1817] ^ m[1818] ^ m[1820] ^ m[1823] ^ m[1825] ^ m[1826] ^ m[1829] ^ m[1830] ^ m[1832] ^ m[1835] ^ m[1836] ^ m[1838] ^ m[1840] ^ m[1843] ^ m[1845] ^ m[1847] ^ m[1848] ^ m[1851] ^ m[1853] ^ m[1854] ^ m[1857] ^ m[1858] ^ m[1860] ^ m[1863] ^ m[1865] ^ m[1866] ^ m[1869] ^ m[1870] ^ m[1872] ^ m[1875] ^ m[1876] ^ m[1878] ^ m[1880] ^ m[1883] ^ m[1885] ^ m[1886] ^ m[1889] ^ m[1890] ^ m[1892] ^ m[1895] ^ m[1896] ^ m[1898] ^ m[1900] ^ m[1903] ^ m[1904] ^ m[1906] ^ m[1908] ^ m[1910] ^ m[1913] ^ m[1915] ^ m[1917] ^ m[1918] ^ m[1921] ^ m[1923] ^ m[1924] ^ m[1927] ^ m[1928] ^ m[1930] ^ m[1933] ^ m[1935] ^ m[1936] ^ m[1939] ^ m[1940] ^ m[1942] ^ m[1945] ^ m[1946] ^ m[1948] ^ m[1950] ^ m[1953] ^ m[1955] ^ m[1956] ^ m[1959] ^ m[1960] ^ m[1962] ^ m[1965] ^ m[1966] ^ m[1968] ^ m[1970] ^ m[1973] ^ m[1974] ^ m[1976] ^ m[1978] ^ m[1980] ^ m[1983] ^ m[1985] ^ m[1986] ^ m[1989] ^ m[1990] ^ m[1992] ^ m[1995] ^ m[1996] ^ m[1998] ^ m[2000] ^ m[2003] ^ m[2004] ^ m[2006] ^ m[2008] ^ m[2010] ^ m[2013] ^ m[2014] ^ m[2016] ^ m[2018] ^ m[2020] ^ m[2022] ^ m[2025] ^ m[2026] ^ m[2027] ^ m[2028] ^ m[2029] ^ m[2030] ^ m[2031] ^ m[2032] ^ m[2033] ^ m[2034] ^ m[2035];
    assign parity[1] = m[1] ^ m[3] ^ m[5] ^ m[7] ^ m[9] ^ m[11] ^ m[13] ^ m[15] ^ m[16] ^ m[19] ^ m[21] ^ m[23] ^ m[25] ^ m[27] ^ m[29] ^ m[31] ^ m[33] ^ m[34] ^ m[37] ^ m[39] ^ m[41] ^ m[43] ^ m[45] ^ m[47] ^ m[49] ^ m[50] ^ m[53] ^ m[55] ^ m[57] ^ m[59] ^ m[61] ^ m[63] ^ m[64] ^ m[67] ^ m[69] ^ m[71] ^ m[73] ^ m[75] ^ m[76] ^ m[79] ^ m[81] ^ m[83] ^ m[85] ^ m[86] ^ m[89] ^ m[91] ^ m[93] ^ m[94] ^ m[97] ^ m[99] ^ m[100] ^ m[103] ^ m[104] ^ m[107] ^ m[108] ^ m[111] ^ m[113] ^ m[115] ^ m[117] ^ m[119] ^ m[121] ^ m[123] ^ m[124] ^ m[127] ^ m[129] ^ m[131] ^ m[133] ^ m[135] ^ m[137] ^ m[139] ^ m[140] ^ m[143] ^ m[145] ^ m[147] ^ m[149] ^ m[151] ^ m[153] ^ m[154] ^ m[157] ^ m[159] ^ m[161] ^ m[163] ^ m[165] ^ m[166] ^ m[169] ^ m[171] ^ m[173] ^ m[175] ^ m[176] ^ m[179] ^ m[181] ^ m[183] ^ m[184] ^ m[187] ^ m[189] ^ m[190] ^ m[193] ^ m[194] ^ m[197] ^ m[198] ^ m[201] ^ m[203] ^ m[205] ^ m[207] ^ m[209] ^ m[211] ^ m[212] ^ m[215] ^ m[217] ^ m[219] ^ m[221] ^ m[223] ^ m[225] ^ m[226] ^ m[229] ^ m[231] ^ m[233] ^ m[235] ^ m[237] ^ m[238] ^ m[241] ^ m[243] ^ m[245] ^ m[247] ^ m[248] ^ m[251] ^ m[253] ^ m[255] ^ m[256] ^ m[259] ^ m[261] ^ m[262] ^ m[265] ^ m[266] ^ m[269] ^ m[270] ^ m[273] ^ m[275] ^ m[277] ^ m[279] ^ m[281] ^ m[282] ^ m[285] ^ m[287] ^ m[289] ^ m[291] ^ m[293] ^ m[294] ^ m[297] ^ m[299] ^ m[301] ^ m[303] ^ m[304] ^ m[307] ^ m[309] ^ m[311] ^ m[312] ^ m[315] ^ m[317] ^ m[318] ^ m[321] ^ m[322] ^ m[325] ^ m[326] ^ m[329] ^ m[331] ^ m[333] ^ m[335] ^ m[336] ^ m[339] ^ m[341] ^ m[343] ^ m[345] ^ m[346] ^ m[349] ^ m[351] ^ m[353] ^ m[354] ^ m[357] ^ m[359] ^ m[360] ^ m[363] ^ m[364] ^ m[367] ^ m[368] ^ m[371] ^ m[373] ^ m[375] ^ m[376] ^ m[379] ^ m[381] ^ m[383] ^ m[384] ^ m[387] ^ m[389] ^ m[390] ^ m[393] ^ m[394] ^ m[397] ^ m[398] ^ m[401] ^ m[403] ^ m[404] ^ m[407] ^ m[409] ^ m[410] ^ m[413] ^ m[414] ^ m[417] ^ m[418] ^ m[421] ^ m[422] ^ m[425] ^ m[426] ^ m[429] ^ m[430] ^ m[432] ^ m[435] ^ m[436] ^ m[438] ^ m[441] ^ m[443] ^ m[445] ^ m[447] ^ m[449] ^ m[451] ^ m[452] ^ m[455] ^ m[457] ^ m[459] ^ m[461] ^ m[463] ^ m[465] ^ m[466] ^ m[469] ^ m[471] ^ m[473] ^ m[475] ^ m[477] ^ m[478] ^ m[481] ^ m[483] ^ m[485] ^ m[487] ^ m[488] ^ m[491] ^ m[493] ^ m[495] ^ m[496] ^ m[499] ^ m[501] ^ m[502] ^ m[505] ^ m[506] ^ m[509] ^ m[510] ^ m[513] ^ m[515] ^ m[517] ^ m[519] ^ m[521] ^ m[522] ^ m[525] ^ m[527] ^ m[529] ^ m[531] ^ m[533] ^ m[534] ^ m[537] ^ m[539] ^ m[541] ^ m[543] ^ m[544] ^ m[547] ^ m[549] ^ m[551] ^ m[552] ^ m[555] ^ m[557] ^ m[558] ^ m[561] ^ m[562] ^ m[565] ^ m[566] ^ m[569] ^ m[571] ^ m[573] ^ m[575] ^ m[576] ^ m[579] ^ m[581] ^ m[583] ^ m[585] ^ m[586] ^ m[589] ^ m[591] ^ m[593] ^ m[594] ^ m[597] ^ m[599] ^ m[600] ^ m[603] ^ m[604] ^ m[607] ^ m[608] ^ m[611] ^ m[613] ^ m[615] ^ m[616] ^ m[619] ^ m[621] ^ m[623] ^ m[624] ^ m[627] ^ m[629] ^ m[630] ^ m[633] ^ m[634] ^ m[637] ^ m[638] ^ m[641] ^ m[643] ^ m[644] ^ m[647] ^ m[649] ^ m[650] ^ m[653] ^ m[654] ^ m[657] ^ m[658] ^ m[661] ^ m[662] ^ m[665] ^ m[666] ^ m[669] ^ m[670] ^ m[672] ^ m[675] ^ m[676] ^ m[678] ^ m[681] ^ m[683] ^ m[685] ^ m[687] ^ m[689] ^ m[690] ^ m[693] ^ m[695] ^ m[697] ^ m[699] ^ m[701] ^ m[702] ^ m[705] ^ m[707] ^ m[709] ^ m[711] ^ m[712] ^ m[715] ^ m[717] ^ m[719] ^ m[720] ^ m[723] ^ m[725] ^ m[726] ^ m[729] ^ m[730] ^ m[733] ^ m[734] ^ m[737] ^ m[739] ^ m[741] ^ m[743] ^ m[744] ^ m[747] ^ m[749] ^ m[751] ^ m[753] ^ m[754] ^ m[757] ^ m[759] ^ m[761] ^ m[762] ^ m[765] ^ m[767] ^ m[768] ^ m[771] ^ m[772] ^ m[775] ^ m[776] ^ m[779] ^ m[781] ^ m[783] ^ m[784] ^ m[787] ^ m[789] ^ m[791] ^ m[792] ^ m[795] ^ m[797] ^ m[798] ^ m[801] ^ m[802] ^ m[805] ^ m[806] ^ m[809] ^ m[811] ^ m[812] ^ m[815] ^ m[817] ^ m[818] ^ m[821] ^ m[822] ^ m[825] ^ m[826] ^ m[829] ^ m[830] ^ m[833] ^ m[834] ^ m[837] ^ m[838] ^ m[840] ^ m[843] ^ m[844] ^ m[846] ^ m[849] ^ m[851] ^ m[853] ^ m[855] ^ m[856] ^ m[859] ^ m[861] ^ m[863] ^ m[865] ^ m[866] ^ m[869] ^ m[871] ^ m[873] ^ m[874] ^ m[877] ^ m[879] ^ m[880] ^ m[883] ^ m[884] ^ m[887] ^ m[888] ^ m[891] ^ m[893] ^ m[895] ^ m[896] ^ m[899] ^ m[901] ^ m[903] ^ m[904] ^ m[907] ^ m[909] ^ m[910] ^ m[913] ^ m[914] ^ m[917] ^ m[918] ^ m[921] ^ m[923] ^ m[924] ^ m[927] ^ m[929] ^ m[930] ^ m[933] ^ m[934] ^ m[937] ^ m[938] ^ m[941] ^ m[942] ^ m[945] ^ m[946] ^ m[949] ^ m[950] ^ m[952] ^ m[955] ^ m[956] ^ m[958] ^ m[961] ^ m[963] ^ m[965] ^ m[966] ^ m[969] ^ m[971] ^ m[973] ^ m[974] ^ m[977] ^ m[979] ^ m[980] ^ m[983] ^ m[984] ^ m[987] ^ m[988] ^ m[991] ^ m[993] ^ m[994] ^ m[997] ^ m[999] ^ m[1000] ^ m[1003] ^ m[1004] ^ m[1007] ^ m[1008] ^ m[1011] ^ m[1012] ^ m[1015] ^ m[1016] ^ m[1019] ^ m[1020] ^ m[1022] ^ m[1025] ^ m[1026] ^ m[1028] ^ m[1031] ^ m[1033] ^ m[1034] ^ m[1037] ^ m[1039] ^ m[1040] ^ m[1043] ^ m[1044] ^ m[1047] ^ m[1048] ^ m[1051] ^ m[1052] ^ m[1055] ^ m[1056] ^ m[1059] ^ m[1060] ^ m[1062] ^ m[1065] ^ m[1066] ^ m[1068] ^ m[1071] ^ m[1072] ^ m[1075] ^ m[1076] ^ m[1079] ^ m[1080] ^ m[1082] ^ m[1085] ^ m[1086] ^ m[1088] ^ m[1090] ^ m[1093] ^ m[1094] ^ m[1096] ^ m[1098] ^ m[1101] ^ m[1103] ^ m[1105] ^ m[1107] ^ m[1109] ^ m[1110] ^ m[1113] ^ m[1115] ^ m[1117] ^ m[1119] ^ m[1121] ^ m[1122] ^ m[1125] ^ m[1127] ^ m[1129] ^ m[1131] ^ m[1132] ^ m[1135] ^ m[1137] ^ m[1139] ^ m[1140] ^ m[1143] ^ m[1145] ^ m[1146] ^ m[1149] ^ m[1150] ^ m[1153] ^ m[1154] ^ m[1157] ^ m[1159] ^ m[1161] ^ m[1163] ^ m[1164] ^ m[1167] ^ m[1169] ^ m[1171] ^ m[1173] ^ m[1174] ^ m[1177] ^ m[1179] ^ m[1181] ^ m[1182] ^ m[1185] ^ m[1187] ^ m[1188] ^ m[1191] ^ m[1192] ^ m[1195] ^ m[1196] ^ m[1199] ^ m[1201] ^ m[1203] ^ m[1204] ^ m[1207] ^ m[1209] ^ m[1211] ^ m[1212] ^ m[1215] ^ m[1217] ^ m[1218] ^ m[1221] ^ m[1222] ^ m[1225] ^ m[1226] ^ m[1229] ^ m[1231] ^ m[1232] ^ m[1235] ^ m[1237] ^ m[1238] ^ m[1241] ^ m[1242] ^ m[1245] ^ m[1246] ^ m[1249] ^ m[1250] ^ m[1253] ^ m[1254] ^ m[1257] ^ m[1258] ^ m[1260] ^ m[1263] ^ m[1264] ^ m[1266] ^ m[1269] ^ m[1271] ^ m[1273] ^ m[1275] ^ m[1276] ^ m[1279] ^ m[1281] ^ m[1283] ^ m[1285] ^ m[1286] ^ m[1289] ^ m[1291] ^ m[1293] ^ m[1294] ^ m[1297] ^ m[1299] ^ m[1300] ^ m[1303] ^ m[1304] ^ m[1307] ^ m[1308] ^ m[1311] ^ m[1313] ^ m[1315] ^ m[1316] ^ m[1319] ^ m[1321] ^ m[1323] ^ m[1324] ^ m[1327] ^ m[1329] ^ m[1330] ^ m[1333] ^ m[1334] ^ m[1337] ^ m[1338] ^ m[1341] ^ m[1343] ^ m[1344] ^ m[1347] ^ m[1349] ^ m[1350] ^ m[1353] ^ m[1354] ^ m[1357] ^ m[1358] ^ m[1361] ^ m[1362] ^ m[1365] ^ m[1366] ^ m[1369] ^ m[1370] ^ m[1372] ^ m[1375] ^ m[1376] ^ m[1378] ^ m[1381] ^ m[1383] ^ m[1385] ^ m[1386] ^ m[1389] ^ m[1391] ^ m[1393] ^ m[1394] ^ m[1397] ^ m[1399] ^ m[1400] ^ m[1403] ^ m[1404] ^ m[1407] ^ m[1408] ^ m[1411] ^ m[1413] ^ m[1414] ^ m[1417] ^ m[1419] ^ m[1420] ^ m[1423] ^ m[1424] ^ m[1427] ^ m[1428] ^ m[1431] ^ m[1432] ^ m[1435] ^ m[1436] ^ m[1439] ^ m[1440] ^ m[1442] ^ m[1445] ^ m[1446] ^ m[1448] ^ m[1451] ^ m[1453] ^ m[1454] ^ m[1457] ^ m[1459] ^ m[1460] ^ m[1463] ^ m[1464] ^ m[1467] ^ m[1468] ^ m[1471] ^ m[1472] ^ m[1475] ^ m[1476] ^ m[1479] ^ m[1480] ^ m[1482] ^ m[1485] ^ m[1486] ^ m[1488] ^ m[1491] ^ m[1492] ^ m[1495] ^ m[1496] ^ m[1499] ^ m[1500] ^ m[1502] ^ m[1505] ^ m[1506] ^ m[1508] ^ m[1510] ^ m[1513] ^ m[1514] ^ m[1516] ^ m[1518] ^ m[1521] ^ m[1523] ^ m[1525] ^ m[1527] ^ m[1528] ^ m[1531] ^ m[1533] ^ m[1535] ^ m[1537] ^ m[1538] ^ m[1541] ^ m[1543] ^ m[1545] ^ m[1546] ^ m[1549] ^ m[1551] ^ m[1552] ^ m[1555] ^ m[1556] ^ m[1559] ^ m[1560] ^ m[1563] ^ m[1565] ^ m[1567] ^ m[1568] ^ m[1571] ^ m[1573] ^ m[1575] ^ m[1576] ^ m[1579] ^ m[1581] ^ m[1582] ^ m[1585] ^ m[1586] ^ m[1589] ^ m[1590] ^ m[1593] ^ m[1595] ^ m[1596] ^ m[1599] ^ m[1601] ^ m[1602] ^ m[1605] ^ m[1606] ^ m[1609] ^ m[1610] ^ m[1613] ^ m[1614] ^ m[1617] ^ m[1618] ^ m[1621] ^ m[1622] ^ m[1624] ^ m[1627] ^ m[1628] ^ m[1630] ^ m[1633] ^ m[1635] ^ m[1637] ^ m[1638] ^ m[1641] ^ m[1643] ^ m[1645] ^ m[1646] ^ m[1649] ^ m[1651] ^ m[1652] ^ m[1655] ^ m[1656] ^ m[1659] ^ m[1660] ^ m[1663] ^ m[1665] ^ m[1666] ^ m[1669] ^ m[1671] ^ m[1672] ^ m[1675] ^ m[1676] ^ m[1679] ^ m[1680] ^ m[1683] ^ m[1684] ^ m[1687] ^ m[1688] ^ m[1691] ^ m[1692] ^ m[1694] ^ m[1697] ^ m[1698] ^ m[1700] ^ m[1703] ^ m[1705] ^ m[1706] ^ m[1709] ^ m[1711] ^ m[1712] ^ m[1715] ^ m[1716] ^ m[1719] ^ m[1720] ^ m[1723] ^ m[1724] ^ m[1727] ^ m[1728] ^ m[1731] ^ m[1732] ^ m[1734] ^ m[1737] ^ m[1738] ^ m[1740] ^ m[1743] ^ m[1744] ^ m[1747] ^ m[1748] ^ m[1751] ^ m[1752] ^ m[1754] ^ m[1757] ^ m[1758] ^ m[1760] ^ m[1762] ^ m[1765] ^ m[1766] ^ m[1768] ^ m[1770] ^ m[1773] ^ m[1775] ^ m[1777] ^ m[1778] ^ m[1781] ^ m[1783] ^ m[1785] ^ m[1786] ^ m[1789] ^ m[1791] ^ m[1792] ^ m[1795] ^ m[1796] ^ m[1799] ^ m[1800] ^ m[1803] ^ m[1805] ^ m[1806] ^ m[1809] ^ m[1811] ^ m[1812] ^ m[1815] ^ m[1816] ^ m[1819] ^ m[1820] ^ m[1823] ^ m[1824] ^ m[1827] ^ m[1828] ^ m[1831] ^ m[1832] ^ m[1834] ^ m[1837] ^ m[1838] ^ m[1840] ^ m[1843] ^ m[1845] ^ m[1846] ^ m[1849] ^ m[1851] ^ m[1852] ^ m[1855] ^ m[1856] ^ m[1859] ^ m[1860] ^ m[1863] ^ m[1864] ^ m[1867] ^ m[1868] ^ m[1871] ^ m[1872] ^ m[1874] ^ m[1877] ^ m[1878] ^ m[1880] ^ m[1883] ^ m[1884] ^ m[1887] ^ m[1888] ^ m[1891] ^ m[1892] ^ m[1894] ^ m[1897] ^ m[1898] ^ m[1900] ^ m[1902] ^ m[1905] ^ m[1906] ^ m[1908] ^ m[1910] ^ m[1913] ^ m[1915] ^ m[1916] ^ m[1919] ^ m[1921] ^ m[1922] ^ m[1925] ^ m[1926] ^ m[1929] ^ m[1930] ^ m[1933] ^ m[1934] ^ m[1937] ^ m[1938] ^ m[1941] ^ m[1942] ^ m[1944] ^ m[1947] ^ m[1948] ^ m[1950] ^ m[1953] ^ m[1954] ^ m[1957] ^ m[1958] ^ m[1961] ^ m[1962] ^ m[1964] ^ m[1967] ^ m[1968] ^ m[1970] ^ m[1972] ^ m[1975] ^ m[1976] ^ m[1978] ^ m[1980] ^ m[1983] ^ m[1984] ^ m[1987] ^ m[1988] ^ m[1991] ^ m[1992] ^ m[1994] ^ m[1997] ^ m[1998] ^ m[2000] ^ m[2002] ^ m[2005] ^ m[2006] ^ m[2008] ^ m[2010] ^ m[2012] ^ m[2015] ^ m[2016] ^ m[2018] ^ m[2020] ^ m[2022] ^ m[2024] ^ m[2026] ^ m[2027] ^ m[2028] ^ m[2029] ^ m[2030] ^ m[2031] ^ m[2032] ^ m[2033] ^ m[2034] ^ m[2035];
    assign parity[2] = m[1] ^ m[3] ^ m[5] ^ m[7] ^ m[9] ^ m[11] ^ m[13] ^ m[14] ^ m[17] ^ m[19] ^ m[21] ^ m[23] ^ m[25] ^ m[27] ^ m[29] ^ m[31] ^ m[32] ^ m[35] ^ m[37] ^ m[39] ^ m[41] ^ m[43] ^ m[45] ^ m[47] ^ m[48] ^ m[51] ^ m[53] ^ m[55] ^ m[57] ^ m[59] ^ m[61] ^ m[62] ^ m[65] ^ m[67] ^ m[69] ^ m[71] ^ m[73] ^ m[74] ^ m[77] ^ m[79] ^ m[81] ^ m[83] ^ m[84] ^ m[87] ^ m[89] ^ m[91] ^ m[92] ^ m[95] ^ m[97] ^ m[98] ^ m[101] ^ m[103] ^ m[104] ^ m[106] ^ m[109] ^ m[111] ^ m[113] ^ m[115] ^ m[117] ^ m[119] ^ m[121] ^ m[122] ^ m[125] ^ m[127] ^ m[129] ^ m[131] ^ m[133] ^ m[135] ^ m[137] ^ m[138] ^ m[141] ^ m[143] ^ m[145] ^ m[147] ^ m[149] ^ m[151] ^ m[152] ^ m[155] ^ m[157] ^ m[159] ^ m[161] ^ m[163] ^ m[164] ^ m[167] ^ m[169] ^ m[171] ^ m[173] ^ m[174] ^ m[177] ^ m[179] ^ m[181] ^ m[182] ^ m[185] ^ m[187] ^ m[188] ^ m[191] ^ m[193] ^ m[194] ^ m[196] ^ m[199] ^ m[201] ^ m[203] ^ m[205] ^ m[207] ^ m[209] ^ m[210] ^ m[213] ^ m[215] ^ m[217] ^ m[219] ^ m[221] ^ m[223] ^ m[224] ^ m[227] ^ m[229] ^ m[231] ^ m[233] ^ m[235] ^ m[236] ^ m[239] ^ m[241] ^ m[243] ^ m[245] ^ m[246] ^ m[249] ^ m[251] ^ m[253] ^ m[254] ^ m[257] ^ m[259] ^ m[260] ^ m[263] ^ m[265] ^ m[266] ^ m[268] ^ m[271] ^ m[273] ^ m[275] ^ m[277] ^ m[279] ^ m[280] ^ m[283] ^ m[285] ^ m[287] ^ m[289] ^ m[291] ^ m[292] ^ m[295] ^ m[297] ^ m[299] ^ m[301] ^ m[302] ^ m[305] ^ m[307] ^ m[309] ^ m[310] ^ m[313] ^ m[315] ^ m[316] ^ m[319] ^ m[321] ^ m[322] ^ m[324] ^ m[327] ^ m[329] ^ m[331] ^ m[333] ^ m[334] ^ m[337] ^ m[339] ^ m[341] ^ m[343] ^ m[344] ^ m[347] ^ m[349] ^ m[351] ^ m[352] ^ m[355] ^ m[357] ^ m[358] ^ m[361] ^ m[363] ^ m[364] ^ m[366] ^ m[369] ^ m[371] ^ m[373] ^ m[374] ^ m[377] ^ m[379] ^ m[381] ^ m[382] ^ m[385] ^ m[387] ^ m[388] ^ m[391] ^ m[393] ^ m[394] ^ m[396] ^ m[399] ^ m[401] ^ m[402] ^ m[405] ^ m[407] ^ m[408] ^ m[411] ^ m[413] ^ m[414] ^ m[416] ^ m[419] ^ m[420] ^ m[423] ^ m[425] ^ m[426] ^ m[428] ^ m[431] ^ m[432] ^ m[434] ^ m[437] ^ m[438] ^ m[441] ^ m[443] ^ m[445] ^ m[447] ^ m[449] ^ m[450] ^ m[453] ^ m[455] ^ m[457] ^ m[459] ^ m[461] ^ m[463] ^ m[464] ^ m[467] ^ m[469] ^ m[471] ^ m[473] ^ m[475] ^ m[476] ^ m[479] ^ m[481] ^ m[483] ^ m[485] ^ m[486] ^ m[489] ^ m[491] ^ m[493] ^ m[494] ^ m[497] ^ m[499] ^ m[500] ^ m[503] ^ m[505] ^ m[506] ^ m[508] ^ m[511] ^ m[513] ^ m[515] ^ m[517] ^ m[519] ^ m[520] ^ m[523] ^ m[525] ^ m[527] ^ m[529] ^ m[531] ^ m[532] ^ m[535] ^ m[537] ^ m[539] ^ m[541] ^ m[542] ^ m[545] ^ m[547] ^ m[549] ^ m[550] ^ m[553] ^ m[555] ^ m[556] ^ m[559] ^ m[561] ^ m[562] ^ m[564] ^ m[567] ^ m[569] ^ m[571] ^ m[573] ^ m[574] ^ m[577] ^ m[579] ^ m[581] ^ m[583] ^ m[584] ^ m[587] ^ m[589] ^ m[591] ^ m[592] ^ m[595] ^ m[597] ^ m[598] ^ m[601] ^ m[603] ^ m[604] ^ m[606] ^ m[609] ^ m[611] ^ m[613] ^ m[614] ^ m[617] ^ m[619] ^ m[621] ^ m[622] ^ m[625] ^ m[627] ^ m[628] ^ m[631] ^ m[633] ^ m[634] ^ m[636] ^ m[639] ^ m[641] ^ m[642] ^ m[645] ^ m[647] ^ m[648] ^ m[651] ^ m[653] ^ m[654] ^ m[656] ^ m[659] ^ m[660] ^ m[663] ^ m[665] ^ m[666] ^ m[668] ^ m[671] ^ m[672] ^ m[674] ^ m[677] ^ m[678] ^ m[681] ^ m[683] ^ m[685] ^ m[687] ^ m[688] ^ m[691] ^ m[693] ^ m[695] ^ m[697] ^ m[699] ^ m[700] ^ m[703] ^ m[705] ^ m[707] ^ m[709] ^ m[710] ^ m[713] ^ m[715] ^ m[717] ^ m[718] ^ m[721] ^ m[723] ^ m[724] ^ m[727] ^ m[729] ^ m[730] ^ m[732] ^ m[735] ^ m[737] ^ m[739] ^ m[741] ^ m[742] ^ m[745] ^ m[747] ^ m[749] ^ m[751] ^ m[752] ^ m[755] ^ m[757] ^ m[759] ^ m[760] ^ m[763] ^ m[765] ^ m[766] ^ m[769] ^ m[771] ^ m[772] ^ m[774] ^ m[777] ^ m[779] ^ m[781] ^ m[782] ^ m[785] ^ m[787] ^ m[789] ^ m[790] ^ m[793] ^ m[795] ^ m[796] ^ m[799] ^ m[801] ^ m[802] ^ m[804] ^ m[807] ^ m[809] ^ m[810] ^ m[813] ^ m[815] ^ m[816] ^ m[819] ^ m[821] ^ m[822] ^ m[824] ^ m[827] ^ m[828] ^ m[831] ^ m[833] ^ m[834] ^ m[836] ^ m[839] ^ m[840] ^ m[842] ^ m[845] ^ m[846] ^ m[849] ^ m[851] ^ m[853] ^ m[854] ^ m[857] ^ m[859] ^ m[861] ^ m[863] ^ m[864] ^ m[867] ^ m[869] ^ m[871] ^ m[872] ^ m[875] ^ m[877] ^ m[878] ^ m[881] ^ m[883] ^ m[884] ^ m[886] ^ m[889] ^ m[891] ^ m[893] ^ m[894] ^ m[897] ^ m[899] ^ m[901] ^ m[902] ^ m[905] ^ m[907] ^ m[908] ^ m[911] ^ m[913] ^ m[914] ^ m[916] ^ m[919] ^ m[921] ^ m[922] ^ m[925] ^ m[927] ^ m[928] ^ m[931] ^ m[933] ^ m[934] ^ m[936] ^ m[939] ^ m[940] ^ m[943] ^ m[945] ^ m[946] ^ m[948] ^ m[951] ^ m[952] ^ m[954] ^ m[957] ^ m[958] ^ m[961] ^ m[963] ^ m[964] ^ m[967] ^ m[969] ^ m[971] ^ m[972] ^ m[975] ^ m[977] ^ m[978] ^ m[981] ^ m[983] ^ m[984] ^ m[986] ^ m[989] ^ m[991] ^ m[992] ^ m[995] ^ m[997] ^ m[998] ^ m[1001] ^ m[1003] ^ m[1004] ^ m[1006] ^ m[1009] ^ m[1010] ^ m[1013] ^ m[1015] ^ m[1016] ^ m[1018] ^ m[1021] ^ m[1022] ^ m[1024] ^ m[1027] ^ m[1028] ^ m[1031] ^ m[1032] ^ m[1035] ^ m[1037] ^ m[1038] ^ m[1041] ^ m[1043] ^ m[1044] ^ m[1046] ^ m[1049] ^ m[1050] ^ m[1053] ^ m[1055] ^ m[1056] ^ m[1058] ^ m[1061] ^ m[1062] ^ m[1064] ^ m[1067] ^ m[1068] ^ m[1070] ^ m[1073] ^ m[1075] ^ m[1076] ^ m[1078] ^ m[1081] ^ m[1082] ^ m[1084] ^ m[1087] ^ m[1088] ^ m[1090] ^ m[1092] ^ m[1095] ^ m[1096] ^ m[1098] ^ m[1101] ^ m[1103] ^ m[1105] ^ m[1107] ^ m[1108] ^ m[1111] ^ m[1113] ^ m[1115] ^ m[1117] ^ m[1119] ^ m[1120] ^ m[1123] ^ m[1125] ^ m[1127] ^ m[1129] ^ m[1130] ^ m[1133] ^ m[1135] ^ m[1137] ^ m[1138] ^ m[1141] ^ m[1143] ^ m[1144] ^ m[1147] ^ m[1149] ^ m[1150] ^ m[1152] ^ m[1155] ^ m[1157] ^ m[1159] ^ m[1161] ^ m[1162] ^ m[1165] ^ m[1167] ^ m[1169] ^ m[1171] ^ m[1172] ^ m[1175] ^ m[1177] ^ m[1179] ^ m[1180] ^ m[1183] ^ m[1185] ^ m[1186] ^ m[1189] ^ m[1191] ^ m[1192] ^ m[1194] ^ m[1197] ^ m[1199] ^ m[1201] ^ m[1202] ^ m[1205] ^ m[1207] ^ m[1209] ^ m[1210] ^ m[1213] ^ m[1215] ^ m[1216] ^ m[1219] ^ m[1221] ^ m[1222] ^ m[1224] ^ m[1227] ^ m[1229] ^ m[1230] ^ m[1233] ^ m[1235] ^ m[1236] ^ m[1239] ^ m[1241] ^ m[1242] ^ m[1244] ^ m[1247] ^ m[1248] ^ m[1251] ^ m[1253] ^ m[1254] ^ m[1256] ^ m[1259] ^ m[1260] ^ m[1262] ^ m[1265] ^ m[1266] ^ m[1269] ^ m[1271] ^ m[1273] ^ m[1274] ^ m[1277] ^ m[1279] ^ m[1281] ^ m[1283] ^ m[1284] ^ m[1287] ^ m[1289] ^ m[1291] ^ m[1292] ^ m[1295] ^ m[1297] ^ m[1298] ^ m[1301] ^ m[1303] ^ m[1304] ^ m[1306] ^ m[1309] ^ m[1311] ^ m[1313] ^ m[1314] ^ m[1317] ^ m[1319] ^ m[1321] ^ m[1322] ^ m[1325] ^ m[1327] ^ m[1328] ^ m[1331] ^ m[1333] ^ m[1334] ^ m[1336] ^ m[1339] ^ m[1341] ^ m[1342] ^ m[1345] ^ m[1347] ^ m[1348] ^ m[1351] ^ m[1353] ^ m[1354] ^ m[1356] ^ m[1359] ^ m[1360] ^ m[1363] ^ m[1365] ^ m[1366] ^ m[1368] ^ m[1371] ^ m[1372] ^ m[1374] ^ m[1377] ^ m[1378] ^ m[1381] ^ m[1383] ^ m[1384] ^ m[1387] ^ m[1389] ^ m[1391] ^ m[1392] ^ m[1395] ^ m[1397] ^ m[1398] ^ m[1401] ^ m[1403] ^ m[1404] ^ m[1406] ^ m[1409] ^ m[1411] ^ m[1412] ^ m[1415] ^ m[1417] ^ m[1418] ^ m[1421] ^ m[1423] ^ m[1424] ^ m[1426] ^ m[1429] ^ m[1430] ^ m[1433] ^ m[1435] ^ m[1436] ^ m[1438] ^ m[1441] ^ m[1442] ^ m[1444] ^ m[1447] ^ m[1448] ^ m[1451] ^ m[1452] ^ m[1455] ^ m[1457] ^ m[1458] ^ m[1461] ^ m[1463] ^ m[1464] ^ m[1466] ^ m[1469] ^ m[1470] ^ m[1473] ^ m[1475] ^ m[1476] ^ m[1478] ^ m[1481] ^ m[1482] ^ m[1484] ^ m[1487] ^ m[1488] ^ m[1490] ^ m[1493] ^ m[1495] ^ m[1496] ^ m[1498] ^ m[1501] ^ m[1502] ^ m[1504] ^ m[1507] ^ m[1508] ^ m[1510] ^ m[1512] ^ m[1515] ^ m[1516] ^ m[1518] ^ m[1521] ^ m[1523] ^ m[1525] ^ m[1526] ^ m[1529] ^ m[1531] ^ m[1533] ^ m[1535] ^ m[1536] ^ m[1539] ^ m[1541] ^ m[1543] ^ m[1544] ^ m[1547] ^ m[1549] ^ m[1550] ^ m[1553] ^ m[1555] ^ m[1556] ^ m[1558] ^ m[1561] ^ m[1563] ^ m[1565] ^ m[1566] ^ m[1569] ^ m[1571] ^ m[1573] ^ m[1574] ^ m[1577] ^ m[1579] ^ m[1580] ^ m[1583] ^ m[1585] ^ m[1586] ^ m[1588] ^ m[1591] ^ m[1593] ^ m[1594] ^ m[1597] ^ m[1599] ^ m[1600] ^ m[1603] ^ m[1605] ^ m[1606] ^ m[1608] ^ m[1611] ^ m[1612] ^ m[1615] ^ m[1617] ^ m[1618] ^ m[1620] ^ m[1623] ^ m[1624] ^ m[1626] ^ m[1629] ^ m[1630] ^ m[1633] ^ m[1635] ^ m[1636] ^ m[1639] ^ m[1641] ^ m[1643] ^ m[1644] ^ m[1647] ^ m[1649] ^ m[1650] ^ m[1653] ^ m[1655] ^ m[1656] ^ m[1658] ^ m[1661] ^ m[1663] ^ m[1664] ^ m[1667] ^ m[1669] ^ m[1670] ^ m[1673] ^ m[1675] ^ m[1676] ^ m[1678] ^ m[1681] ^ m[1682] ^ m[1685] ^ m[1687] ^ m[1688] ^ m[1690] ^ m[1693] ^ m[1694] ^ m[1696] ^ m[1699] ^ m[1700] ^ m[1703] ^ m[1704] ^ m[1707] ^ m[1709] ^ m[1710] ^ m[1713] ^ m[1715] ^ m[1716] ^ m[1718] ^ m[1721] ^ m[1722] ^ m[1725] ^ m[1727] ^ m[1728] ^ m[1730] ^ m[1733] ^ m[1734] ^ m[1736] ^ m[1739] ^ m[1740] ^ m[1742] ^ m[1745] ^ m[1747] ^ m[1748] ^ m[1750] ^ m[1753] ^ m[1754] ^ m[1756] ^ m[1759] ^ m[1760] ^ m[1762] ^ m[1764] ^ m[1767] ^ m[1768] ^ m[1770] ^ m[1773] ^ m[1775] ^ m[1776] ^ m[1779] ^ m[1781] ^ m[1783] ^ m[1784] ^ m[1787] ^ m[1789] ^ m[1790] ^ m[1793] ^ m[1795] ^ m[1796] ^ m[1798] ^ m[1801] ^ m[1803] ^ m[1804] ^ m[1807] ^ m[1809] ^ m[1810] ^ m[1813] ^ m[1815] ^ m[1816] ^ m[1818] ^ m[1821] ^ m[1822] ^ m[1825] ^ m[1827] ^ m[1828] ^ m[1830] ^ m[1833] ^ m[1834] ^ m[1836] ^ m[1839] ^ m[1840] ^ m[1843] ^ m[1844] ^ m[1847] ^ m[1849] ^ m[1850] ^ m[1853] ^ m[1855] ^ m[1856] ^ m[1858] ^ m[1861] ^ m[1862] ^ m[1865] ^ m[1867] ^ m[1868] ^ m[1870] ^ m[1873] ^ m[1874] ^ m[1876] ^ m[1879] ^ m[1880] ^ m[1882] ^ m[1885] ^ m[1887] ^ m[1888] ^ m[1890] ^ m[1893] ^ m[1894] ^ m[1896] ^ m[1899] ^ m[1900] ^ m[1902] ^ m[1904] ^ m[1907] ^ m[1908] ^ m[1910] ^ m[1913] ^ m[1914] ^ m[1917] ^ m[1919] ^ m[1920] ^ m[1923] ^ m[1925] ^ m[1926] ^ m[1928] ^ m[1931] ^ m[1932] ^ m[1935] ^ m[1937] ^ m[1938] ^ m[1940] ^ m[1943] ^ m[1944] ^ m[1946] ^ m[1949] ^ m[1950] ^ m[1952] ^ m[1955] ^ m[1957] ^ m[1958] ^ m[1960] ^ m[1963] ^ m[1964] ^ m[1966] ^ m[1969] ^ m[1970] ^ m[1972] ^ m[1974] ^ m[1977] ^ m[1978] ^ m[1980] ^ m[1982] ^ m[1985] ^ m[1987] ^ m[1988] ^ m[1990] ^ m[1993] ^ m[1994] ^ m[1996] ^ m[1999] ^ m[2000] ^ m[2002] ^ m[2004] ^ m[2007] ^ m[2008] ^ m[2010] ^ m[2012] ^ m[2014] ^ m[2017] ^ m[2018] ^ m[2020] ^ m[2022] ^ m[2024] ^ m[2025] ^ m[2027] ^ m[2028] ^ m[2029] ^ m[2030] ^ m[2031] ^ m[2032] ^ m[2033] ^ m[2034] ^ m[2035];
    assign parity[3] = m[1] ^ m[3] ^ m[5] ^ m[7] ^ m[9] ^ m[11] ^ m[12] ^ m[15] ^ m[17] ^ m[19] ^ m[21] ^ m[23] ^ m[25] ^ m[27] ^ m[29] ^ m[30] ^ m[33] ^ m[35] ^ m[37] ^ m[39] ^ m[41] ^ m[43] ^ m[45] ^ m[46] ^ m[49] ^ m[51] ^ m[53] ^ m[55] ^ m[57] ^ m[59] ^ m[60] ^ m[63] ^ m[65] ^ m[67] ^ m[69] ^ m[71] ^ m[72] ^ m[75] ^ m[77] ^ m[79] ^ m[81] ^ m[82] ^ m[85] ^ m[87] ^ m[89] ^ m[90] ^ m[93] ^ m[95] ^ m[97] ^ m[98] ^ m[100] ^ m[102] ^ m[105] ^ m[107] ^ m[109] ^ m[111] ^ m[113] ^ m[115] ^ m[117] ^ m[119] ^ m[120] ^ m[123] ^ m[125] ^ m[127] ^ m[129] ^ m[131] ^ m[133] ^ m[135] ^ m[136] ^ m[139] ^ m[141] ^ m[143] ^ m[145] ^ m[147] ^ m[149] ^ m[150] ^ m[153] ^ m[155] ^ m[157] ^ m[159] ^ m[161] ^ m[162] ^ m[165] ^ m[167] ^ m[169] ^ m[171] ^ m[172] ^ m[175] ^ m[177] ^ m[179] ^ m[180] ^ m[183] ^ m[185] ^ m[187] ^ m[188] ^ m[190] ^ m[192] ^ m[195] ^ m[197] ^ m[199] ^ m[201] ^ m[203] ^ m[205] ^ m[207] ^ m[208] ^ m[211] ^ m[213] ^ m[215] ^ m[217] ^ m[219] ^ m[221] ^ m[222] ^ m[225] ^ m[227] ^ m[229] ^ m[231] ^ m[233] ^ m[234] ^ m[237] ^ m[239] ^ m[241] ^ m[243] ^ m[244] ^ m[247] ^ m[249] ^ m[251] ^ m[252] ^ m[255] ^ m[257] ^ m[259] ^ m[260] ^ m[262] ^ m[264] ^ m[267] ^ m[269] ^ m[271] ^ m[273] ^ m[275] ^ m[277] ^ m[278] ^ m[281] ^ m[283] ^ m[285] ^ m[287] ^ m[289] ^ m[290] ^ m[293] ^ m[295] ^ m[297] ^ m[299] ^ m[300] ^ m[303] ^ m[305] ^ m[307] ^ m[308] ^ m[311] ^ m[313] ^ m[315] ^ m[316] ^ m[318] ^ m[320] ^ m[323] ^ m[325] ^ m[327] ^ m[329] ^ m[331] ^ m[332] ^ m[335] ^ m[337] ^ m[339] ^ m[341] ^ m[342] ^ m[345] ^ m[347] ^ m[349] ^ m[350] ^ m[353] ^ m[355] ^ m[357] ^ m[358] ^ m[360] ^ m[362] ^ m[365] ^ m[367] ^ m[369] ^ m[371] ^ m[372] ^ m[375] ^ m[377] ^ m[379] ^ m[380] ^ m[383] ^ m[385] ^ m[387] ^ m[388] ^ m[390] ^ m[392] ^ m[395] ^ m[397] ^ m[399] ^ m[400] ^ m[403] ^ m[405] ^ m[407] ^ m[408] ^ m[410] ^ m[412] ^ m[415] ^ m[417] ^ m[419] ^ m[420] ^ m[422] ^ m[424] ^ m[427] ^ m[429] ^ m[431] ^ m[432] ^ m[434] ^ m[436] ^ m[439] ^ m[441] ^ m[443] ^ m[445] ^ m[447] ^ m[448] ^ m[451] ^ m[453] ^ m[455] ^ m[457] ^ m[459] ^ m[461] ^ m[462] ^ m[465] ^ m[467] ^ m[469] ^ m[471] ^ m[473] ^ m[474] ^ m[477] ^ m[479] ^ m[481] ^ m[483] ^ m[484] ^ m[487] ^ m[489] ^ m[491] ^ m[492] ^ m[495] ^ m[497] ^ m[499] ^ m[500] ^ m[502] ^ m[504] ^ m[507] ^ m[509] ^ m[511] ^ m[513] ^ m[515] ^ m[517] ^ m[518] ^ m[521] ^ m[523] ^ m[525] ^ m[527] ^ m[529] ^ m[530] ^ m[533] ^ m[535] ^ m[537] ^ m[539] ^ m[540] ^ m[543] ^ m[545] ^ m[547] ^ m[548] ^ m[551] ^ m[553] ^ m[555] ^ m[556] ^ m[558] ^ m[560] ^ m[563] ^ m[565] ^ m[567] ^ m[569] ^ m[571] ^ m[572] ^ m[575] ^ m[577] ^ m[579] ^ m[581] ^ m[582] ^ m[585] ^ m[587] ^ m[589] ^ m[590] ^ m[593] ^ m[595] ^ m[597] ^ m[598] ^ m[600] ^ m[602] ^ m[605] ^ m[607] ^ m[609] ^ m[611] ^ m[612] ^ m[615] ^ m[617] ^ m[619] ^ m[620] ^ m[623] ^ m[625] ^ m[627] ^ m[628] ^ m[630] ^ m[632] ^ m[635] ^ m[637] ^ m[639] ^ m[640] ^ m[643] ^ m[645] ^ m[647] ^ m[648] ^ m[650] ^ m[652] ^ m[655] ^ m[657] ^ m[659] ^ m[660] ^ m[662] ^ m[664] ^ m[667] ^ m[669] ^ m[671] ^ m[672] ^ m[674] ^ m[676] ^ m[679] ^ m[681] ^ m[683] ^ m[685] ^ m[686] ^ m[689] ^ m[691] ^ m[693] ^ m[695] ^ m[697] ^ m[698] ^ m[701] ^ m[703] ^ m[705] ^ m[707] ^ m[708] ^ m[711] ^ m[713] ^ m[715] ^ m[716] ^ m[719] ^ m[721] ^ m[723] ^ m[724] ^ m[726] ^ m[728] ^ m[731] ^ m[733] ^ m[735] ^ m[737] ^ m[739] ^ m[740] ^ m[743] ^ m[745] ^ m[747] ^ m[749] ^ m[750] ^ m[753] ^ m[755] ^ m[757] ^ m[758] ^ m[761] ^ m[763] ^ m[765] ^ m[766] ^ m[768] ^ m[770] ^ m[773] ^ m[775] ^ m[777] ^ m[779] ^ m[780] ^ m[783] ^ m[785] ^ m[787] ^ m[788] ^ m[791] ^ m[793] ^ m[795] ^ m[796] ^ m[798] ^ m[800] ^ m[803] ^ m[805] ^ m[807] ^ m[808] ^ m[811] ^ m[813] ^ m[815] ^ m[816] ^ m[818] ^ m[820] ^ m[823] ^ m[825] ^ m[827] ^ m[828] ^ m[830] ^ m[832] ^ m[835] ^ m[837] ^ m[839] ^ m[840] ^ m[842] ^ m[844] ^ m[847] ^ m[849] ^ m[851] ^ m[852] ^ m[855] ^ m[857] ^ m[859] ^ m[861] ^ m[862] ^ m[865] ^ m[867] ^ m[869] ^ m[870] ^ m[873] ^ m[875] ^ m[877] ^ m[878] ^ m[880] ^ m[882] ^ m[885] ^ m[887] ^ m[889] ^ m[891] ^ m[892] ^ m[895] ^ m[897] ^ m[899] ^ m[900] ^ m[903] ^ m[905] ^ m[907] ^ m[908] ^ m[910] ^ m[912] ^ m[915] ^ m[917] ^ m[919] ^ m[920] ^ m[923] ^ m[925] ^ m[927] ^ m[928] ^ m[930] ^ m[932] ^ m[935] ^ m[937] ^ m[939] ^ m[940] ^ m[942] ^ m[944] ^ m[947] ^ m[949] ^ m[951] ^ m[952] ^ m[954] ^ m[956] ^ m[959] ^ m[961] ^ m[962] ^ m[965] ^ m[967] ^ m[969] ^ m[970] ^ m[973] ^ m[975] ^ m[977] ^ m[978] ^ m[980] ^ m[982] ^ m[985] ^ m[987] ^ m[989] ^ m[990] ^ m[993] ^ m[995] ^ m[997] ^ m[998] ^ m[1000] ^ m[1002] ^ m[1005] ^ m[1007] ^ m[1009] ^ m[1010] ^ m[1012] ^ m[1014] ^ m[1017] ^ m[1019] ^ m[1021] ^ m[1022] ^ m[1024] ^ m[1026] ^ m[1029] ^ m[1030] ^ m[1033] ^ m[1035] ^ m[1037] ^ m[1038] ^ m[1040] ^ m[1042] ^ m[1045] ^ m[1047] ^ m[1049] ^ m[1050] ^ m[1052] ^ m[1054] ^ m[1057] ^ m[1059] ^ m[1061] ^ m[1062] ^ m[1064] ^ m[1066] ^ m[1069] ^ m[1070] ^ m[1072] ^ m[1074] ^ m[1077] ^ m[1079] ^ m[1081] ^ m[1082] ^ m[1084] ^ m[1086] ^ m[1089] ^ m[1090] ^ m[1092] ^ m[1094] ^ m[1097] ^ m[1098] ^ m[1101] ^ m[1103] ^ m[1105] ^ m[1106] ^ m[1109] ^ m[1111] ^ m[1113] ^ m[1115] ^ m[1117] ^ m[1118] ^ m[1121] ^ m[1123] ^ m[1125] ^ m[1127] ^ m[1128] ^ m[1131] ^ m[1133] ^ m[1135] ^ m[1136] ^ m[1139] ^ m[1141] ^ m[1143] ^ m[1144] ^ m[1146] ^ m[1148] ^ m[1151] ^ m[1153] ^ m[1155] ^ m[1157] ^ m[1159] ^ m[1160] ^ m[1163] ^ m[1165] ^ m[1167] ^ m[1169] ^ m[1170] ^ m[1173] ^ m[1175] ^ m[1177] ^ m[1178] ^ m[1181] ^ m[1183] ^ m[1185] ^ m[1186] ^ m[1188] ^ m[1190] ^ m[1193] ^ m[1195] ^ m[1197] ^ m[1199] ^ m[1200] ^ m[1203] ^ m[1205] ^ m[1207] ^ m[1208] ^ m[1211] ^ m[1213] ^ m[1215] ^ m[1216] ^ m[1218] ^ m[1220] ^ m[1223] ^ m[1225] ^ m[1227] ^ m[1228] ^ m[1231] ^ m[1233] ^ m[1235] ^ m[1236] ^ m[1238] ^ m[1240] ^ m[1243] ^ m[1245] ^ m[1247] ^ m[1248] ^ m[1250] ^ m[1252] ^ m[1255] ^ m[1257] ^ m[1259] ^ m[1260] ^ m[1262] ^ m[1264] ^ m[1267] ^ m[1269] ^ m[1271] ^ m[1272] ^ m[1275] ^ m[1277] ^ m[1279] ^ m[1281] ^ m[1282] ^ m[1285] ^ m[1287] ^ m[1289] ^ m[1290] ^ m[1293] ^ m[1295] ^ m[1297] ^ m[1298] ^ m[1300] ^ m[1302] ^ m[1305] ^ m[1307] ^ m[1309] ^ m[1311] ^ m[1312] ^ m[1315] ^ m[1317] ^ m[1319] ^ m[1320] ^ m[1323] ^ m[1325] ^ m[1327] ^ m[1328] ^ m[1330] ^ m[1332] ^ m[1335] ^ m[1337] ^ m[1339] ^ m[1340] ^ m[1343] ^ m[1345] ^ m[1347] ^ m[1348] ^ m[1350] ^ m[1352] ^ m[1355] ^ m[1357] ^ m[1359] ^ m[1360] ^ m[1362] ^ m[1364] ^ m[1367] ^ m[1369] ^ m[1371] ^ m[1372] ^ m[1374] ^ m[1376] ^ m[1379] ^ m[1381] ^ m[1382] ^ m[1385] ^ m[1387] ^ m[1389] ^ m[1390] ^ m[1393] ^ m[1395] ^ m[1397] ^ m[1398] ^ m[1400] ^ m[1402] ^ m[1405] ^ m[1407] ^ m[1409] ^ m[1410] ^ m[1413] ^ m[1415] ^ m[1417] ^ m[1418] ^ m[1420] ^ m[1422] ^ m[1425] ^ m[1427] ^ m[1429] ^ m[1430] ^ m[1432] ^ m[1434] ^ m[1437] ^ m[1439] ^ m[1441] ^ m[1442] ^ m[1444] ^ m[1446] ^ m[1449] ^ m[1450] ^ m[1453] ^ m[1455] ^ m[1457] ^ m[1458] ^ m[1460] ^ m[1462] ^ m[1465] ^ m[1467] ^ m[1469] ^ m[1470] ^ m[1472] ^ m[1474] ^ m[1477] ^ m[1479] ^ m[1481] ^ m[1482] ^ m[1484] ^ m[1486] ^ m[1489] ^ m[1490] ^ m[1492] ^ m[1494] ^ m[1497] ^ m[1499] ^ m[1501] ^ m[1502] ^ m[1504] ^ m[1506] ^ m[1509] ^ m[1510] ^ m[1512] ^ m[1514] ^ m[1517] ^ m[1518] ^ m[1521] ^ m[1523] ^ m[1524] ^ m[1527] ^ m[1529] ^ m[1531] ^ m[1533] ^ m[1534] ^ m[1537] ^ m[1539] ^ m[1541] ^ m[1542] ^ m[1545] ^ m[1547] ^ m[1549] ^ m[1550] ^ m[1552] ^ m[1554] ^ m[1557] ^ m[1559] ^ m[1561] ^ m[1563] ^ m[1564] ^ m[1567] ^ m[1569] ^ m[1571] ^ m[1572] ^ m[1575] ^ m[1577] ^ m[1579] ^ m[1580] ^ m[1582] ^ m[1584] ^ m[1587] ^ m[1589] ^ m[1591] ^ m[1592] ^ m[1595] ^ m[1597] ^ m[1599] ^ m[1600] ^ m[1602] ^ m[1604] ^ m[1607] ^ m[1609] ^ m[1611] ^ m[1612] ^ m[1614] ^ m[1616] ^ m[1619] ^ m[1621] ^ m[1623] ^ m[1624] ^ m[1626] ^ m[1628] ^ m[1631] ^ m[1633] ^ m[1634] ^ m[1637] ^ m[1639] ^ m[1641] ^ m[1642] ^ m[1645] ^ m[1647] ^ m[1649] ^ m[1650] ^ m[1652] ^ m[1654] ^ m[1657] ^ m[1659] ^ m[1661] ^ m[1662] ^ m[1665] ^ m[1667] ^ m[1669] ^ m[1670] ^ m[1672] ^ m[1674] ^ m[1677] ^ m[1679] ^ m[1681] ^ m[1682] ^ m[1684] ^ m[1686] ^ m[1689] ^ m[1691] ^ m[1693] ^ m[1694] ^ m[1696] ^ m[1698] ^ m[1701] ^ m[1702] ^ m[1705] ^ m[1707] ^ m[1709] ^ m[1710] ^ m[1712] ^ m[1714] ^ m[1717] ^ m[1719] ^ m[1721] ^ m[1722] ^ m[1724] ^ m[1726] ^ m[1729] ^ m[1731] ^ m[1733] ^ m[1734] ^ m[1736] ^ m[1738] ^ m[1741] ^ m[1742] ^ m[1744] ^ m[1746] ^ m[1749] ^ m[1751] ^ m[1753] ^ m[1754] ^ m[1756] ^ m[1758] ^ m[1761] ^ m[1762] ^ m[1764] ^ m[1766] ^ m[1769] ^ m[1770] ^ m[1773] ^ m[1774] ^ m[1777] ^ m[1779] ^ m[1781] ^ m[1782] ^ m[1785] ^ m[1787] ^ m[1789] ^ m[1790] ^ m[1792] ^ m[1794] ^ m[1797] ^ m[1799] ^ m[1801] ^ m[1802] ^ m[1805] ^ m[1807] ^ m[1809] ^ m[1810] ^ m[1812] ^ m[1814] ^ m[1817] ^ m[1819] ^ m[1821] ^ m[1822] ^ m[1824] ^ m[1826] ^ m[1829] ^ m[1831] ^ m[1833] ^ m[1834] ^ m[1836] ^ m[1838] ^ m[1841] ^ m[1842] ^ m[1845] ^ m[1847] ^ m[1849] ^ m[1850] ^ m[1852] ^ m[1854] ^ m[1857] ^ m[1859] ^ m[1861] ^ m[1862] ^ m[1864] ^ m[1866] ^ m[1869] ^ m[1871] ^ m[1873] ^ m[1874] ^ m[1876] ^ m[1878] ^ m[1881] ^ m[1882] ^ m[1884] ^ m[1886] ^ m[1889] ^ m[1891] ^ m[1893] ^ m[1894] ^ m[1896] ^ m[1898] ^ m[1901] ^ m[1902] ^ m[1904] ^ m[1906] ^ m[1909] ^ m[1910] ^ m[1912] ^ m[1915] ^ m[1917] ^ m[1919] ^ m[1920] ^ m[1922] ^ m[1924] ^ m[1927] ^ m[1929] ^ m[1931] ^ m[1932] ^ m[1934] ^ m[1936] ^ m[1939] ^ m[1941] ^ m[1943] ^ m[1944] ^ m[1946] ^ m[1948] ^ m[1951] ^ m[1952] ^ m[1954] ^ m[1956] ^ m[1959] ^ m[1961] ^ m[1963] ^ m[1964] ^ m[1966] ^ m[1968] ^ m[1971] ^ m[1972] ^ m[1974] ^ m[1976] ^ m[1979] ^ m[1980] ^ m[1982] ^ m[1984] ^ m[1986] ^ m[1989] ^ m[1991] ^ m[1993] ^ m[1994] ^ m[1996] ^ m[1998] ^ m[2001] ^ m[2002] ^ m[2004] ^ m[2006] ^ m[2009] ^ m[2010] ^ m[2012] ^ m[2014] ^ m[2016] ^ m[2019] ^ m[2020] ^ m[2022] ^ m[2024] ^ m[2025] ^ m[2026] ^ m[2028] ^ m[2029] ^ m[2030] ^ m[2031] ^ m[2032] ^ m[2033] ^ m[2034] ^ m[2035];
    assign parity[4] = m[1] ^ m[3] ^ m[5] ^ m[7] ^ m[9] ^ m[10] ^ m[13] ^ m[15] ^ m[17] ^ m[19] ^ m[21] ^ m[23] ^ m[25] ^ m[27] ^ m[28] ^ m[31] ^ m[33] ^ m[35] ^ m[37] ^ m[39] ^ m[41] ^ m[43] ^ m[44] ^ m[47] ^ m[49] ^ m[51] ^ m[53] ^ m[55] ^ m[57] ^ m[58] ^ m[61] ^ m[63] ^ m[65] ^ m[67] ^ m[69] ^ m[70] ^ m[73] ^ m[75] ^ m[77] ^ m[79] ^ m[80] ^ m[83] ^ m[85] ^ m[87] ^ m[89] ^ m[90] ^ m[92] ^ m[94] ^ m[96] ^ m[99] ^ m[101] ^ m[103] ^ m[105] ^ m[107] ^ m[109] ^ m[111] ^ m[113] ^ m[115] ^ m[117] ^ m[118] ^ m[121] ^ m[123] ^ m[125] ^ m[127] ^ m[129] ^ m[131] ^ m[133] ^ m[134] ^ m[137] ^ m[139] ^ m[141] ^ m[143] ^ m[145] ^ m[147] ^ m[148] ^ m[151] ^ m[153] ^ m[155] ^ m[157] ^ m[159] ^ m[160] ^ m[163] ^ m[165] ^ m[167] ^ m[169] ^ m[170] ^ m[173] ^ m[175] ^ m[177] ^ m[179] ^ m[180] ^ m[182] ^ m[184] ^ m[186] ^ m[189] ^ m[191] ^ m[193] ^ m[195] ^ m[197] ^ m[199] ^ m[201] ^ m[203] ^ m[205] ^ m[206] ^ m[209] ^ m[211] ^ m[213] ^ m[215] ^ m[217] ^ m[219] ^ m[220] ^ m[223] ^ m[225] ^ m[227] ^ m[229] ^ m[231] ^ m[232] ^ m[235] ^ m[237] ^ m[239] ^ m[241] ^ m[242] ^ m[245] ^ m[247] ^ m[249] ^ m[251] ^ m[252] ^ m[254] ^ m[256] ^ m[258] ^ m[261] ^ m[263] ^ m[265] ^ m[267] ^ m[269] ^ m[271] ^ m[273] ^ m[275] ^ m[276] ^ m[279] ^ m[281] ^ m[283] ^ m[285] ^ m[287] ^ m[288] ^ m[291] ^ m[293] ^ m[295] ^ m[297] ^ m[298] ^ m[301] ^ m[303] ^ m[305] ^ m[307] ^ m[308] ^ m[310] ^ m[312] ^ m[314] ^ m[317] ^ m[319] ^ m[321] ^ m[323] ^ m[325] ^ m[327] ^ m[329] ^ m[330] ^ m[333] ^ m[335] ^ m[337] ^ m[339] ^ m[340] ^ m[343] ^ m[345] ^ m[347] ^ m[349] ^ m[350] ^ m[352] ^ m[354] ^ m[356] ^ m[359] ^ m[361] ^ m[363] ^ m[365] ^ m[367] ^ m[369] ^ m[370] ^ m[373] ^ m[375] ^ m[377] ^ m[379] ^ m[380] ^ m[382] ^ m[384] ^ m[386] ^ m[389] ^ m[391] ^ m[393] ^ m[395] ^ m[397] ^ m[399] ^ m[400] ^ m[402] ^ m[404] ^ m[406] ^ m[409] ^ m[411] ^ m[413] ^ m[415] ^ m[417] ^ m[419] ^ m[420] ^ m[422] ^ m[424] ^ m[426] ^ m[428] ^ m[430] ^ m[433] ^ m[435] ^ m[437] ^ m[439] ^ m[441] ^ m[443] ^ m[445] ^ m[446] ^ m[449] ^ m[451] ^ m[453] ^ m[455] ^ m[457] ^ m[459] ^ m[460] ^ m[463] ^ m[465] ^ m[467] ^ m[469] ^ m[471] ^ m[472] ^ m[475] ^ m[477] ^ m[479] ^ m[481] ^ m[482] ^ m[485] ^ m[487] ^ m[489] ^ m[491] ^ m[492] ^ m[494] ^ m[496] ^ m[498] ^ m[501] ^ m[503] ^ m[505] ^ m[507] ^ m[509] ^ m[511] ^ m[513] ^ m[515] ^ m[516] ^ m[519] ^ m[521] ^ m[523] ^ m[525] ^ m[527] ^ m[528] ^ m[531] ^ m[533] ^ m[535] ^ m[537] ^ m[538] ^ m[541] ^ m[543] ^ m[545] ^ m[547] ^ m[548] ^ m[550] ^ m[552] ^ m[554] ^ m[557] ^ m[559] ^ m[561] ^ m[563] ^ m[565] ^ m[567] ^ m[569] ^ m[570] ^ m[573] ^ m[575] ^ m[577] ^ m[579] ^ m[580] ^ m[583] ^ m[585] ^ m[587] ^ m[589] ^ m[590] ^ m[592] ^ m[594] ^ m[596] ^ m[599] ^ m[601] ^ m[603] ^ m[605] ^ m[607] ^ m[609] ^ m[610] ^ m[613] ^ m[615] ^ m[617] ^ m[619] ^ m[620] ^ m[622] ^ m[624] ^ m[626] ^ m[629] ^ m[631] ^ m[633] ^ m[635] ^ m[637] ^ m[639] ^ m[640] ^ m[642] ^ m[644] ^ m[646] ^ m[649] ^ m[651] ^ m[653] ^ m[655] ^ m[657] ^ m[659] ^ m[660] ^ m[662] ^ m[664] ^ m[666] ^ m[668] ^ m[670] ^ m[673] ^ m[675] ^ m[677] ^ m[679] ^ m[681] ^ m[683] ^ m[684] ^ m[687] ^ m[689] ^ m[691] ^ m[693] ^ m[695] ^ m[696] ^ m[699] ^ m[701] ^ m[703] ^ m[705] ^ m[706] ^ m[709] ^ m[711] ^ m[713] ^ m[715] ^ m[716] ^ m[718] ^ m[720] ^ m[722] ^ m[725] ^ m[727] ^ m[729] ^ m[731] ^ m[733] ^ m[735] ^ m[737] ^ m[738] ^ m[741] ^ m[743] ^ m[745] ^ m[747] ^ m[748] ^ m[751] ^ m[753] ^ m[755] ^ m[757] ^ m[758] ^ m[760] ^ m[762] ^ m[764] ^ m[767] ^ m[769] ^ m[771] ^ m[773] ^ m[775] ^ m[777] ^ m[778] ^ m[781] ^ m[783] ^ m[785] ^ m[787] ^ m[788] ^ m[790] ^ m[792] ^ m[794] ^ m[797] ^ m[799] ^ m[801] ^ m[803] ^ m[805] ^ m[807] ^ m[808] ^ m[810] ^ m[812] ^ m[814] ^ m[817] ^ m[819] ^ m[821] ^ m[823] ^ m[825] ^ m[827] ^ m[828] ^ m[830] ^ m[832] ^ m[834] ^ m[836] ^ m[838] ^ m[841] ^ m[843] ^ m[845] ^ m[847] ^ m[849] ^ m[850] ^ m[853] ^ m[855] ^ m[857] ^ m[859] ^ m[860] ^ m[863] ^ m[865] ^ m[867] ^ m[869] ^ m[870] ^ m[872] ^ m[874] ^ m[876] ^ m[879] ^ m[881] ^ m[883] ^ m[885] ^ m[887] ^ m[889] ^ m[890] ^ m[893] ^ m[895] ^ m[897] ^ m[899] ^ m[900] ^ m[902] ^ m[904] ^ m[906] ^ m[909] ^ m[911] ^ m[913] ^ m[915] ^ m[917] ^ m[919] ^ m[920] ^ m[922] ^ m[924] ^ m[926] ^ m[929] ^ m[931] ^ m[933] ^ m[935] ^ m[937] ^ m[939] ^ m[940] ^ m[942] ^ m[944] ^ m[946] ^ m[948] ^ m[950] ^ m[953] ^ m[955] ^ m[957] ^ m[959] ^ m[960] ^ m[963] ^ m[965] ^ m[967] ^ m[969] ^ m[970] ^ m[972] ^ m[974] ^ m[976] ^ m[979] ^ m[981] ^ m[983] ^ m[985] ^ m[987] ^ m[989] ^ m[990] ^ m[992] ^ m[994] ^ m[996] ^ m[999] ^ m[1001] ^ m[1003] ^ m[1005] ^ m[1007] ^ m[1009] ^ m[1010] ^ m[1012] ^ m[1014] ^ m[1016] ^ m[1018] ^ m[1020] ^ m[1023] ^ m[1025] ^ m[1027] ^ m[1029] ^ m[1030] ^ m[1032] ^ m[1034] ^ m[1036] ^ m[1039] ^ m[1041] ^ m[1043] ^ m[1045] ^ m[1047] ^ m[1049] ^ m[1050] ^ m[1052] ^ m[1054] ^ m[1056] ^ m[1058] ^ m[1060] ^ m[1063] ^ m[1065] ^ m[1067] ^ m[1069] ^ m[1070] ^ m[1072] ^ m[1074] ^ m[1076] ^ m[1078] ^ m[1080] ^ m[1083] ^ m[1085] ^ m[1087] ^ m[1089] ^ m[1090] ^ m[1092] ^ m[1094] ^ m[1096] ^ m[1099] ^ m[1101] ^ m[1103] ^ m[1104] ^ m[1107] ^ m[1109] ^ m[1111] ^ m[1113] ^ m[1115] ^ m[1116] ^ m[1119] ^ m[1121] ^ m[1123] ^ m[1125] ^ m[1126] ^ m[1129] ^ m[1131] ^ m[1133] ^ m[1135] ^ m[1136] ^ m[1138] ^ m[1140] ^ m[1142] ^ m[1145] ^ m[1147] ^ m[1149] ^ m[1151] ^ m[1153] ^ m[1155] ^ m[1157] ^ m[1158] ^ m[1161] ^ m[1163] ^ m[1165] ^ m[1167] ^ m[1168] ^ m[1171] ^ m[1173] ^ m[1175] ^ m[1177] ^ m[1178] ^ m[1180] ^ m[1182] ^ m[1184] ^ m[1187] ^ m[1189] ^ m[1191] ^ m[1193] ^ m[1195] ^ m[1197] ^ m[1198] ^ m[1201] ^ m[1203] ^ m[1205] ^ m[1207] ^ m[1208] ^ m[1210] ^ m[1212] ^ m[1214] ^ m[1217] ^ m[1219] ^ m[1221] ^ m[1223] ^ m[1225] ^ m[1227] ^ m[1228] ^ m[1230] ^ m[1232] ^ m[1234] ^ m[1237] ^ m[1239] ^ m[1241] ^ m[1243] ^ m[1245] ^ m[1247] ^ m[1248] ^ m[1250] ^ m[1252] ^ m[1254] ^ m[1256] ^ m[1258] ^ m[1261] ^ m[1263] ^ m[1265] ^ m[1267] ^ m[1269] ^ m[1270] ^ m[1273] ^ m[1275] ^ m[1277] ^ m[1279] ^ m[1280] ^ m[1283] ^ m[1285] ^ m[1287] ^ m[1289] ^ m[1290] ^ m[1292] ^ m[1294] ^ m[1296] ^ m[1299] ^ m[1301] ^ m[1303] ^ m[1305] ^ m[1307] ^ m[1309] ^ m[1310] ^ m[1313] ^ m[1315] ^ m[1317] ^ m[1319] ^ m[1320] ^ m[1322] ^ m[1324] ^ m[1326] ^ m[1329] ^ m[1331] ^ m[1333] ^ m[1335] ^ m[1337] ^ m[1339] ^ m[1340] ^ m[1342] ^ m[1344] ^ m[1346] ^ m[1349] ^ m[1351] ^ m[1353] ^ m[1355] ^ m[1357] ^ m[1359] ^ m[1360] ^ m[1362] ^ m[1364] ^ m[1366] ^ m[1368] ^ m[1370] ^ m[1373] ^ m[1375] ^ m[1377] ^ m[1379] ^ m[1380] ^ m[1383] ^ m[1385] ^ m[1387] ^ m[1389] ^ m[1390] ^ m[1392] ^ m[1394] ^ m[1396] ^ m[1399] ^ m[1401] ^ m[1403] ^ m[1405] ^ m[1407] ^ m[1409] ^ m[1410] ^ m[1412] ^ m[1414] ^ m[1416] ^ m[1419] ^ m[1421] ^ m[1423] ^ m[1425] ^ m[1427] ^ m[1429] ^ m[1430] ^ m[1432] ^ m[1434] ^ m[1436] ^ m[1438] ^ m[1440] ^ m[1443] ^ m[1445] ^ m[1447] ^ m[1449] ^ m[1450] ^ m[1452] ^ m[1454] ^ m[1456] ^ m[1459] ^ m[1461] ^ m[1463] ^ m[1465] ^ m[1467] ^ m[1469] ^ m[1470] ^ m[1472] ^ m[1474] ^ m[1476] ^ m[1478] ^ m[1480] ^ m[1483] ^ m[1485] ^ m[1487] ^ m[1489] ^ m[1490] ^ m[1492] ^ m[1494] ^ m[1496] ^ m[1498] ^ m[1500] ^ m[1503] ^ m[1505] ^ m[1507] ^ m[1509] ^ m[1510] ^ m[1512] ^ m[1514] ^ m[1516] ^ m[1519] ^ m[1521] ^ m[1522] ^ m[1525] ^ m[1527] ^ m[1529] ^ m[1531] ^ m[1532] ^ m[1535] ^ m[1537] ^ m[1539] ^ m[1541] ^ m[1542] ^ m[1544] ^ m[1546] ^ m[1548] ^ m[1551] ^ m[1553] ^ m[1555] ^ m[1557] ^ m[1559] ^ m[1561] ^ m[1562] ^ m[1565] ^ m[1567] ^ m[1569] ^ m[1571] ^ m[1572] ^ m[1574] ^ m[1576] ^ m[1578] ^ m[1581] ^ m[1583] ^ m[1585] ^ m[1587] ^ m[1589] ^ m[1591] ^ m[1592] ^ m[1594] ^ m[1596] ^ m[1598] ^ m[1601] ^ m[1603] ^ m[1605] ^ m[1607] ^ m[1609] ^ m[1611] ^ m[1612] ^ m[1614] ^ m[1616] ^ m[1618] ^ m[1620] ^ m[1622] ^ m[1625] ^ m[1627] ^ m[1629] ^ m[1631] ^ m[1632] ^ m[1635] ^ m[1637] ^ m[1639] ^ m[1641] ^ m[1642] ^ m[1644] ^ m[1646] ^ m[1648] ^ m[1651] ^ m[1653] ^ m[1655] ^ m[1657] ^ m[1659] ^ m[1661] ^ m[1662] ^ m[1664] ^ m[1666] ^ m[1668] ^ m[1671] ^ m[1673] ^ m[1675] ^ m[1677] ^ m[1679] ^ m[1681] ^ m[1682] ^ m[1684] ^ m[1686] ^ m[1688] ^ m[1690] ^ m[1692] ^ m[1695] ^ m[1697] ^ m[1699] ^ m[1701] ^ m[1702] ^ m[1704] ^ m[1706] ^ m[1708] ^ m[1711] ^ m[1713] ^ m[1715] ^ m[1717] ^ m[1719] ^ m[1721] ^ m[1722] ^ m[1724] ^ m[1726] ^ m[1728] ^ m[1730] ^ m[1732] ^ m[1735] ^ m[1737] ^ m[1739] ^ m[1741] ^ m[1742] ^ m[1744] ^ m[1746] ^ m[1748] ^ m[1750] ^ m[1752] ^ m[1755] ^ m[1757] ^ m[1759] ^ m[1761] ^ m[1762] ^ m[1764] ^ m[1766] ^ m[1768] ^ m[1771] ^ m[1772] ^ m[1775] ^ m[1777] ^ m[1779] ^ m[1781] ^ m[1782] ^ m[1784] ^ m[1786] ^ m[1788] ^ m[1791] ^ m[1793] ^ m[1795] ^ m[1797] ^ m[1799] ^ m[1801] ^ m[1802] ^ m[1804] ^ m[1806] ^ m[1808] ^ m[1811] ^ m[1813] ^ m[1815] ^ m[1817] ^ m[1819] ^ m[1821] ^ m[1822] ^ m[1824] ^ m[1826] ^ m[1828] ^ m[1830] ^ m[1832] ^ m[1835] ^ m[1837] ^ m[1839] ^ m[1841] ^ m[1842] ^ m[1844] ^ m[1846] ^ m[1848] ^ m[1851] ^ m[1853] ^ m[1855] ^ m[1857] ^ m[1859] ^ m[1861] ^ m[1862] ^ m[1864] ^ m[1866] ^ m[1868] ^ m[1870] ^ m[1872] ^ m[1875] ^ m[1877] ^ m[1879] ^ m[1881] ^ m[1882] ^ m[1884] ^ m[1886] ^ m[1888] ^ m[1890] ^ m[1892] ^ m[1895] ^ m[1897] ^ m[1899] ^ m[1901] ^ m[1902] ^ m[1904] ^ m[1906] ^ m[1908] ^ m[1911] ^ m[1912] ^ m[1914] ^ m[1916] ^ m[1918] ^ m[1921] ^ m[1923] ^ m[1925] ^ m[1927] ^ m[1929] ^ m[1931] ^ m[1932] ^ m[1934] ^ m[1936] ^ m[1938] ^ m[1940] ^ m[1942] ^ m[1945] ^ m[1947] ^ m[1949] ^ m[1951] ^ m[1952] ^ m[1954] ^ m[1956] ^ m[1958] ^ m[1960] ^ m[1962] ^ m[1965] ^ m[1967] ^ m[1969] ^ m[1971] ^ m[1972] ^ m[1974] ^ m[1976] ^ m[1978] ^ m[1981] ^ m[1982] ^ m[1984] ^ m[1986] ^ m[1988] ^ m[1990] ^ m[1992] ^ m[1995] ^ m[1997] ^ m[1999] ^ m[2001] ^ m[2002] ^ m[2004] ^ m[2006] ^ m[2008] ^ m[2011] ^ m[2012] ^ m[2014] ^ m[2016] ^ m[2018] ^ m[2021] ^ m[2022] ^ m[2024] ^ m[2025] ^ m[2026] ^ m[2027] ^ m[2029] ^ m[2030] ^ m[2031] ^ m[2032] ^ m[2033] ^ m[2034] ^ m[2035];
    assign parity[5] = m[1] ^ m[3] ^ m[5] ^ m[7] ^ m[8] ^ m[11] ^ m[13] ^ m[15] ^ m[17] ^ m[19] ^ m[21] ^ m[23] ^ m[25] ^ m[26] ^ m[29] ^ m[31] ^ m[33] ^ m[35] ^ m[37] ^ m[39] ^ m[41] ^ m[42] ^ m[45] ^ m[47] ^ m[49] ^ m[51] ^ m[53] ^ m[55] ^ m[56] ^ m[59] ^ m[61] ^ m[63] ^ m[65] ^ m[67] ^ m[68] ^ m[71] ^ m[73] ^ m[75] ^ m[77] ^ m[79] ^ m[80] ^ m[82] ^ m[84] ^ m[86] ^ m[88] ^ m[91] ^ m[93] ^ m[95] ^ m[97] ^ m[99] ^ m[101] ^ m[103] ^ m[105] ^ m[107] ^ m[109] ^ m[111] ^ m[113] ^ m[115] ^ m[116] ^ m[119] ^ m[121] ^ m[123] ^ m[125] ^ m[127] ^ m[129] ^ m[131] ^ m[132] ^ m[135] ^ m[137] ^ m[139] ^ m[141] ^ m[143] ^ m[145] ^ m[146] ^ m[149] ^ m[151] ^ m[153] ^ m[155] ^ m[157] ^ m[158] ^ m[161] ^ m[163] ^ m[165] ^ m[167] ^ m[169] ^ m[170] ^ m[172] ^ m[174] ^ m[176] ^ m[178] ^ m[181] ^ m[183] ^ m[185] ^ m[187] ^ m[189] ^ m[191] ^ m[193] ^ m[195] ^ m[197] ^ m[199] ^ m[201] ^ m[203] ^ m[204] ^ m[207] ^ m[209] ^ m[211] ^ m[213] ^ m[215] ^ m[217] ^ m[218] ^ m[221] ^ m[223] ^ m[225] ^ m[227] ^ m[229] ^ m[230] ^ m[233] ^ m[235] ^ m[237] ^ m[239] ^ m[241] ^ m[242] ^ m[244] ^ m[246] ^ m[248] ^ m[250] ^ m[253] ^ m[255] ^ m[257] ^ m[259] ^ m[261] ^ m[263] ^ m[265] ^ m[267] ^ m[269] ^ m[271] ^ m[273] ^ m[274] ^ m[277] ^ m[279] ^ m[281] ^ m[283] ^ m[285] ^ m[286] ^ m[289] ^ m[291] ^ m[293] ^ m[295] ^ m[297] ^ m[298] ^ m[300] ^ m[302] ^ m[304] ^ m[306] ^ m[309] ^ m[311] ^ m[313] ^ m[315] ^ m[317] ^ m[319] ^ m[321] ^ m[323] ^ m[325] ^ m[327] ^ m[328] ^ m[331] ^ m[333] ^ m[335] ^ m[337] ^ m[339] ^ m[340] ^ m[342] ^ m[344] ^ m[346] ^ m[348] ^ m[351] ^ m[353] ^ m[355] ^ m[357] ^ m[359] ^ m[361] ^ m[363] ^ m[365] ^ m[367] ^ m[369] ^ m[370] ^ m[372] ^ m[374] ^ m[376] ^ m[378] ^ m[381] ^ m[383] ^ m[385] ^ m[387] ^ m[389] ^ m[391] ^ m[393] ^ m[395] ^ m[397] ^ m[399] ^ m[400] ^ m[402] ^ m[404] ^ m[406] ^ m[408] ^ m[410] ^ m[412] ^ m[414] ^ m[416] ^ m[418] ^ m[421] ^ m[423] ^ m[425] ^ m[427] ^ m[429] ^ m[431] ^ m[433] ^ m[435] ^ m[437] ^ m[439] ^ m[441] ^ m[443] ^ m[444] ^ m[447] ^ m[449] ^ m[451] ^ m[453] ^ m[455] ^ m[457] ^ m[458] ^ m[461] ^ m[463] ^ m[465] ^ m[467] ^ m[469] ^ m[470] ^ m[473] ^ m[475] ^ m[477] ^ m[479] ^ m[481] ^ m[482] ^ m[484] ^ m[486] ^ m[488] ^ m[490] ^ m[493] ^ m[495] ^ m[497] ^ m[499] ^ m[501] ^ m[503] ^ m[505] ^ m[507] ^ m[509] ^ m[511] ^ m[513] ^ m[514] ^ m[517] ^ m[519] ^ m[521] ^ m[523] ^ m[525] ^ m[526] ^ m[529] ^ m[531] ^ m[533] ^ m[535] ^ m[537] ^ m[538] ^ m[540] ^ m[542] ^ m[544] ^ m[546] ^ m[549] ^ m[551] ^ m[553] ^ m[555] ^ m[557] ^ m[559] ^ m[561] ^ m[563] ^ m[565] ^ m[567] ^ m[568] ^ m[571] ^ m[573] ^ m[575] ^ m[577] ^ m[579] ^ m[580] ^ m[582] ^ m[584] ^ m[586] ^ m[588] ^ m[591] ^ m[593] ^ m[595] ^ m[597] ^ m[599] ^ m[601] ^ m[603] ^ m[605] ^ m[607] ^ m[609] ^ m[610] ^ m[612] ^ m[614] ^ m[616] ^ m[618] ^ m[621] ^ m[623] ^ m[625] ^ m[627] ^ m[629] ^ m[631] ^ m[633] ^ m[635] ^ m[637] ^ m[639] ^ m[640] ^ m[642] ^ m[644] ^ m[646] ^ m[648] ^ m[650] ^ m[652] ^ m[654] ^ m[656] ^ m[658] ^ m[661] ^ m[663] ^ m[665] ^ m[667] ^ m[669] ^ m[671] ^ m[673] ^ m[675] ^ m[677] ^ m[679] ^ m[681] ^ m[682] ^ m[685] ^ m[687] ^ m[689] ^ m[691] ^ m[693] ^ m[694] ^ m[697] ^ m[699] ^ m[701] ^ m[703] ^ m[705] ^ m[706] ^ m[708] ^ m[710] ^ m[712] ^ m[714] ^ m[717] ^ m[719] ^ m[721] ^ m[723] ^ m[725] ^ m[727] ^ m[729] ^ m[731] ^ m[733] ^ m[735] ^ m[736] ^ m[739] ^ m[741] ^ m[743] ^ m[745] ^ m[747] ^ m[748] ^ m[750] ^ m[752] ^ m[754] ^ m[756] ^ m[759] ^ m[761] ^ m[763] ^ m[765] ^ m[767] ^ m[769] ^ m[771] ^ m[773] ^ m[775] ^ m[777] ^ m[778] ^ m[780] ^ m[782] ^ m[784] ^ m[786] ^ m[789] ^ m[791] ^ m[793] ^ m[795] ^ m[797] ^ m[799] ^ m[801] ^ m[803] ^ m[805] ^ m[807] ^ m[808] ^ m[810] ^ m[812] ^ m[814] ^ m[816] ^ m[818] ^ m[820] ^ m[822] ^ m[824] ^ m[826] ^ m[829] ^ m[831] ^ m[833] ^ m[835] ^ m[837] ^ m[839] ^ m[841] ^ m[843] ^ m[845] ^ m[847] ^ m[848] ^ m[851] ^ m[853] ^ m[855] ^ m[857] ^ m[859] ^ m[860] ^ m[862] ^ m[864] ^ m[866] ^ m[868] ^ m[871] ^ m[873] ^ m[875] ^ m[877] ^ m[879] ^ m[881] ^ m[883] ^ m[885] ^ m[887] ^ m[889] ^ m[890] ^ m[892] ^ m[894] ^ m[896] ^ m[898] ^ m[901] ^ m[903] ^ m[905] ^ m[907] ^ m[909] ^ m[911] ^ m[913] ^ m[915] ^ m[917] ^ m[919] ^ m[920] ^ m[922] ^ m[924] ^ m[926] ^ m[928] ^ m[930] ^ m[932] ^ m[934] ^ m[936] ^ m[938] ^ m[941] ^ m[943] ^ m[945] ^ m[947] ^ m[949] ^ m[951] ^ m[953] ^ m[955] ^ m[957] ^ m[959] ^ m[960] ^ m[962] ^ m[964] ^ m[966] ^ m[968] ^ m[971] ^ m[973] ^ m[975] ^ m[977] ^ m[979] ^ m[981] ^ m[983] ^ m[985] ^ m[987] ^ m[989] ^ m[990] ^ m[992] ^ m[994] ^ m[996] ^ m[998] ^ m[1000] ^ m[1002] ^ m[1004] ^ m[1006] ^ m[1008] ^ m[1011] ^ m[1013] ^ m[1015] ^ m[1017] ^ m[1019] ^ m[1021] ^ m[1023] ^ m[1025] ^ m[1027] ^ m[1029] ^ m[1030] ^ m[1032] ^ m[1034] ^ m[1036] ^ m[1038] ^ m[1040] ^ m[1042] ^ m[1044] ^ m[1046] ^ m[1048] ^ m[1051] ^ m[1053] ^ m[1055] ^ m[1057] ^ m[1059] ^ m[1061] ^ m[1063] ^ m[1065] ^ m[1067] ^ m[1069] ^ m[1070] ^ m[1072] ^ m[1074] ^ m[1076] ^ m[1078] ^ m[1080] ^ m[1082] ^ m[1084] ^ m[1086] ^ m[1088] ^ m[1091] ^ m[1093] ^ m[1095] ^ m[1097] ^ m[1099] ^ m[1101] ^ m[1102] ^ m[1105] ^ m[1107] ^ m[1109] ^ m[1111] ^ m[1113] ^ m[1114] ^ m[1117] ^ m[1119] ^ m[1121] ^ m[1123] ^ m[1125] ^ m[1126] ^ m[1128] ^ m[1130] ^ m[1132] ^ m[1134] ^ m[1137] ^ m[1139] ^ m[1141] ^ m[1143] ^ m[1145] ^ m[1147] ^ m[1149] ^ m[1151] ^ m[1153] ^ m[1155] ^ m[1156] ^ m[1159] ^ m[1161] ^ m[1163] ^ m[1165] ^ m[1167] ^ m[1168] ^ m[1170] ^ m[1172] ^ m[1174] ^ m[1176] ^ m[1179] ^ m[1181] ^ m[1183] ^ m[1185] ^ m[1187] ^ m[1189] ^ m[1191] ^ m[1193] ^ m[1195] ^ m[1197] ^ m[1198] ^ m[1200] ^ m[1202] ^ m[1204] ^ m[1206] ^ m[1209] ^ m[1211] ^ m[1213] ^ m[1215] ^ m[1217] ^ m[1219] ^ m[1221] ^ m[1223] ^ m[1225] ^ m[1227] ^ m[1228] ^ m[1230] ^ m[1232] ^ m[1234] ^ m[1236] ^ m[1238] ^ m[1240] ^ m[1242] ^ m[1244] ^ m[1246] ^ m[1249] ^ m[1251] ^ m[1253] ^ m[1255] ^ m[1257] ^ m[1259] ^ m[1261] ^ m[1263] ^ m[1265] ^ m[1267] ^ m[1268] ^ m[1271] ^ m[1273] ^ m[1275] ^ m[1277] ^ m[1279] ^ m[1280] ^ m[1282] ^ m[1284] ^ m[1286] ^ m[1288] ^ m[1291] ^ m[1293] ^ m[1295] ^ m[1297] ^ m[1299] ^ m[1301] ^ m[1303] ^ m[1305] ^ m[1307] ^ m[1309] ^ m[1310] ^ m[1312] ^ m[1314] ^ m[1316] ^ m[1318] ^ m[1321] ^ m[1323] ^ m[1325] ^ m[1327] ^ m[1329] ^ m[1331] ^ m[1333] ^ m[1335] ^ m[1337] ^ m[1339] ^ m[1340] ^ m[1342] ^ m[1344] ^ m[1346] ^ m[1348] ^ m[1350] ^ m[1352] ^ m[1354] ^ m[1356] ^ m[1358] ^ m[1361] ^ m[1363] ^ m[1365] ^ m[1367] ^ m[1369] ^ m[1371] ^ m[1373] ^ m[1375] ^ m[1377] ^ m[1379] ^ m[1380] ^ m[1382] ^ m[1384] ^ m[1386] ^ m[1388] ^ m[1391] ^ m[1393] ^ m[1395] ^ m[1397] ^ m[1399] ^ m[1401] ^ m[1403] ^ m[1405] ^ m[1407] ^ m[1409] ^ m[1410] ^ m[1412] ^ m[1414] ^ m[1416] ^ m[1418] ^ m[1420] ^ m[1422] ^ m[1424] ^ m[1426] ^ m[1428] ^ m[1431] ^ m[1433] ^ m[1435] ^ m[1437] ^ m[1439] ^ m[1441] ^ m[1443] ^ m[1445] ^ m[1447] ^ m[1449] ^ m[1450] ^ m[1452] ^ m[1454] ^ m[1456] ^ m[1458] ^ m[1460] ^ m[1462] ^ m[1464] ^ m[1466] ^ m[1468] ^ m[1471] ^ m[1473] ^ m[1475] ^ m[1477] ^ m[1479] ^ m[1481] ^ m[1483] ^ m[1485] ^ m[1487] ^ m[1489] ^ m[1490] ^ m[1492] ^ m[1494] ^ m[1496] ^ m[1498] ^ m[1500] ^ m[1502] ^ m[1504] ^ m[1506] ^ m[1508] ^ m[1511] ^ m[1513] ^ m[1515] ^ m[1517] ^ m[1519] ^ m[1520] ^ m[1523] ^ m[1525] ^ m[1527] ^ m[1529] ^ m[1531] ^ m[1532] ^ m[1534] ^ m[1536] ^ m[1538] ^ m[1540] ^ m[1543] ^ m[1545] ^ m[1547] ^ m[1549] ^ m[1551] ^ m[1553] ^ m[1555] ^ m[1557] ^ m[1559] ^ m[1561] ^ m[1562] ^ m[1564] ^ m[1566] ^ m[1568] ^ m[1570] ^ m[1573] ^ m[1575] ^ m[1577] ^ m[1579] ^ m[1581] ^ m[1583] ^ m[1585] ^ m[1587] ^ m[1589] ^ m[1591] ^ m[1592] ^ m[1594] ^ m[1596] ^ m[1598] ^ m[1600] ^ m[1602] ^ m[1604] ^ m[1606] ^ m[1608] ^ m[1610] ^ m[1613] ^ m[1615] ^ m[1617] ^ m[1619] ^ m[1621] ^ m[1623] ^ m[1625] ^ m[1627] ^ m[1629] ^ m[1631] ^ m[1632] ^ m[1634] ^ m[1636] ^ m[1638] ^ m[1640] ^ m[1643] ^ m[1645] ^ m[1647] ^ m[1649] ^ m[1651] ^ m[1653] ^ m[1655] ^ m[1657] ^ m[1659] ^ m[1661] ^ m[1662] ^ m[1664] ^ m[1666] ^ m[1668] ^ m[1670] ^ m[1672] ^ m[1674] ^ m[1676] ^ m[1678] ^ m[1680] ^ m[1683] ^ m[1685] ^ m[1687] ^ m[1689] ^ m[1691] ^ m[1693] ^ m[1695] ^ m[1697] ^ m[1699] ^ m[1701] ^ m[1702] ^ m[1704] ^ m[1706] ^ m[1708] ^ m[1710] ^ m[1712] ^ m[1714] ^ m[1716] ^ m[1718] ^ m[1720] ^ m[1723] ^ m[1725] ^ m[1727] ^ m[1729] ^ m[1731] ^ m[1733] ^ m[1735] ^ m[1737] ^ m[1739] ^ m[1741] ^ m[1742] ^ m[1744] ^ m[1746] ^ m[1748] ^ m[1750] ^ m[1752] ^ m[1754] ^ m[1756] ^ m[1758] ^ m[1760] ^ m[1763] ^ m[1765] ^ m[1767] ^ m[1769] ^ m[1771] ^ m[1772] ^ m[1774] ^ m[1776] ^ m[1778] ^ m[1780] ^ m[1783] ^ m[1785] ^ m[1787] ^ m[1789] ^ m[1791] ^ m[1793] ^ m[1795] ^ m[1797] ^ m[1799] ^ m[1801] ^ m[1802] ^ m[1804] ^ m[1806] ^ m[1808] ^ m[1810] ^ m[1812] ^ m[1814] ^ m[1816] ^ m[1818] ^ m[1820] ^ m[1823] ^ m[1825] ^ m[1827] ^ m[1829] ^ m[1831] ^ m[1833] ^ m[1835] ^ m[1837] ^ m[1839] ^ m[1841] ^ m[1842] ^ m[1844] ^ m[1846] ^ m[1848] ^ m[1850] ^ m[1852] ^ m[1854] ^ m[1856] ^ m[1858] ^ m[1860] ^ m[1863] ^ m[1865] ^ m[1867] ^ m[1869] ^ m[1871] ^ m[1873] ^ m[1875] ^ m[1877] ^ m[1879] ^ m[1881] ^ m[1882] ^ m[1884] ^ m[1886] ^ m[1888] ^ m[1890] ^ m[1892] ^ m[1894] ^ m[1896] ^ m[1898] ^ m[1900] ^ m[1903] ^ m[1905] ^ m[1907] ^ m[1909] ^ m[1911] ^ m[1912] ^ m[1914] ^ m[1916] ^ m[1918] ^ m[1920] ^ m[1922] ^ m[1924] ^ m[1926] ^ m[1928] ^ m[1930] ^ m[1933] ^ m[1935] ^ m[1937] ^ m[1939] ^ m[1941] ^ m[1943] ^ m[1945] ^ m[1947] ^ m[1949] ^ m[1951] ^ m[1952] ^ m[1954] ^ m[1956] ^ m[1958] ^ m[1960] ^ m[1962] ^ m[1964] ^ m[1966] ^ m[1968] ^ m[1970] ^ m[1973] ^ m[1975] ^ m[1977] ^ m[1979] ^ m[1981] ^ m[1982] ^ m[1984] ^ m[1986] ^ m[1988] ^ m[1990] ^ m[1992] ^ m[1994] ^ m[1996] ^ m[1998] ^ m[2000] ^ m[2003] ^ m[2005] ^ m[2007] ^ m[2009] ^ m[2011] ^ m[2012] ^ m[2014] ^ m[2016] ^ m[2018] ^ m[2020] ^ m[2023] ^ m[2024] ^ m[2025] ^ m[2026] ^ m[2027] ^ m[2028] ^ m[2030] ^ m[2031] ^ m[2032] ^ m[2033] ^ m[2034] ^ m[2035];
    assign parity[6] = m[1] ^ m[3] ^ m[5] ^ m[6] ^ m[9] ^ m[11] ^ m[13] ^ m[15] ^ m[17] ^ m[19] ^ m[21] ^ m[23] ^ m[24] ^ m[27] ^ m[29] ^ m[31] ^ m[33] ^ m[35] ^ m[37] ^ m[39] ^ m[40] ^ m[43] ^ m[45] ^ m[47] ^ m[49] ^ m[51] ^ m[53] ^ m[54] ^ m[57] ^ m[59] ^ m[61] ^ m[63] ^ m[65] ^ m[67] ^ m[68] ^ m[70] ^ m[72] ^ m[74] ^ m[76] ^ m[78] ^ m[81] ^ m[83] ^ m[85] ^ m[87] ^ m[89] ^ m[91] ^ m[93] ^ m[95] ^ m[97] ^ m[99] ^ m[101] ^ m[103] ^ m[105] ^ m[107] ^ m[109] ^ m[111] ^ m[113] ^ m[114] ^ m[117] ^ m[119] ^ m[121] ^ m[123] ^ m[125] ^ m[127] ^ m[129] ^ m[130] ^ m[133] ^ m[135] ^ m[137] ^ m[139] ^ m[141] ^ m[143] ^ m[144] ^ m[147] ^ m[149] ^ m[151] ^ m[153] ^ m[155] ^ m[157] ^ m[158] ^ m[160] ^ m[162] ^ m[164] ^ m[166] ^ m[168] ^ m[171] ^ m[173] ^ m[175] ^ m[177] ^ m[179] ^ m[181] ^ m[183] ^ m[185] ^ m[187] ^ m[189] ^ m[191] ^ m[193] ^ m[195] ^ m[197] ^ m[199] ^ m[201] ^ m[202] ^ m[205] ^ m[207] ^ m[209] ^ m[211] ^ m[213] ^ m[215] ^ m[216] ^ m[219] ^ m[221] ^ m[223] ^ m[225] ^ m[227] ^ m[229] ^ m[230] ^ m[232] ^ m[234] ^ m[236] ^ m[238] ^ m[240] ^ m[243] ^ m[245] ^ m[247] ^ m[249] ^ m[251] ^ m[253] ^ m[255] ^ m[257] ^ m[259] ^ m[261] ^ m[263] ^ m[265] ^ m[267] ^ m[269] ^ m[271] ^ m[272] ^ m[275] ^ m[277] ^ m[279] ^ m[281] ^ m[283] ^ m[285] ^ m[286] ^ m[288] ^ m[290] ^ m[292] ^ m[294] ^ m[296] ^ m[299] ^ m[301] ^ m[303] ^ m[305] ^ m[307] ^ m[309] ^ m[311] ^ m[313] ^ m[315] ^ m[317] ^ m[319] ^ m[321] ^ m[323] ^ m[325] ^ m[327] ^ m[328] ^ m[330] ^ m[332] ^ m[334] ^ m[336] ^ m[338] ^ m[341] ^ m[343] ^ m[345] ^ m[347] ^ m[349] ^ m[351] ^ m[353] ^ m[355] ^ m[357] ^ m[359] ^ m[361] ^ m[363] ^ m[365] ^ m[367] ^ m[369] ^ m[370] ^ m[372] ^ m[374] ^ m[376] ^ m[378] ^ m[380] ^ m[382] ^ m[384] ^ m[386] ^ m[388] ^ m[390] ^ m[392] ^ m[394] ^ m[396] ^ m[398] ^ m[401] ^ m[403] ^ m[405] ^ m[407] ^ m[409] ^ m[411] ^ m[413] ^ m[415] ^ m[417] ^ m[419] ^ m[421] ^ m[423] ^ m[425] ^ m[427] ^ m[429] ^ m[431] ^ m[433] ^ m[435] ^ m[437] ^ m[439] ^ m[441] ^ m[442] ^ m[445] ^ m[447] ^ m[449] ^ m[451] ^ m[453] ^ m[455] ^ m[456] ^ m[459] ^ m[461] ^ m[463] ^ m[465] ^ m[467] ^ m[469] ^ m[470] ^ m[472] ^ m[474] ^ m[476] ^ m[478] ^ m[480] ^ m[483] ^ m[485] ^ m[487] ^ m[489] ^ m[491] ^ m[493] ^ m[495] ^ m[497] ^ m[499] ^ m[501] ^ m[503] ^ m[505] ^ m[507] ^ m[509] ^ m[511] ^ m[512] ^ m[515] ^ m[517] ^ m[519] ^ m[521] ^ m[523] ^ m[525] ^ m[526] ^ m[528] ^ m[530] ^ m[532] ^ m[534] ^ m[536] ^ m[539] ^ m[541] ^ m[543] ^ m[545] ^ m[547] ^ m[549] ^ m[551] ^ m[553] ^ m[555] ^ m[557] ^ m[559] ^ m[561] ^ m[563] ^ m[565] ^ m[567] ^ m[568] ^ m[570] ^ m[572] ^ m[574] ^ m[576] ^ m[578] ^ m[581] ^ m[583] ^ m[585] ^ m[587] ^ m[589] ^ m[591] ^ m[593] ^ m[595] ^ m[597] ^ m[599] ^ m[601] ^ m[603] ^ m[605] ^ m[607] ^ m[609] ^ m[610] ^ m[612] ^ m[614] ^ m[616] ^ m[618] ^ m[620] ^ m[622] ^ m[624] ^ m[626] ^ m[628] ^ m[630] ^ m[632] ^ m[634] ^ m[636] ^ m[638] ^ m[641] ^ m[643] ^ m[645] ^ m[647] ^ m[649] ^ m[651] ^ m[653] ^ m[655] ^ m[657] ^ m[659] ^ m[661] ^ m[663] ^ m[665] ^ m[667] ^ m[669] ^ m[671] ^ m[673] ^ m[675] ^ m[677] ^ m[679] ^ m[680] ^ m[683] ^ m[685] ^ m[687] ^ m[689] ^ m[691] ^ m[693] ^ m[694] ^ m[696] ^ m[698] ^ m[700] ^ m[702] ^ m[704] ^ m[707] ^ m[709] ^ m[711] ^ m[713] ^ m[715] ^ m[717] ^ m[719] ^ m[721] ^ m[723] ^ m[725] ^ m[727] ^ m[729] ^ m[731] ^ m[733] ^ m[735] ^ m[736] ^ m[738] ^ m[740] ^ m[742] ^ m[744] ^ m[746] ^ m[749] ^ m[751] ^ m[753] ^ m[755] ^ m[757] ^ m[759] ^ m[761] ^ m[763] ^ m[765] ^ m[767] ^ m[769] ^ m[771] ^ m[773] ^ m[775] ^ m[777] ^ m[778] ^ m[780] ^ m[782] ^ m[784] ^ m[786] ^ m[788] ^ m[790] ^ m[792] ^ m[794] ^ m[796] ^ m[798] ^ m[800] ^ m[802] ^ m[804] ^ m[806] ^ m[809] ^ m[811] ^ m[813] ^ m[815] ^ m[817] ^ m[819] ^ m[821] ^ m[823] ^ m[825] ^ m[827] ^ m[829] ^ m[831] ^ m[833] ^ m[835] ^ m[837] ^ m[839] ^ m[841] ^ m[843] ^ m[845] ^ m[847] ^ m[848] ^ m[850] ^ m[852] ^ m[854] ^ m[856] ^ m[858] ^ m[861] ^ m[863] ^ m[865] ^ m[867] ^ m[869] ^ m[871] ^ m[873] ^ m[875] ^ m[877] ^ m[879] ^ m[881] ^ m[883] ^ m[885] ^ m[887] ^ m[889] ^ m[890] ^ m[892] ^ m[894] ^ m[896] ^ m[898] ^ m[900] ^ m[902] ^ m[904] ^ m[906] ^ m[908] ^ m[910] ^ m[912] ^ m[914] ^ m[916] ^ m[918] ^ m[921] ^ m[923] ^ m[925] ^ m[927] ^ m[929] ^ m[931] ^ m[933] ^ m[935] ^ m[937] ^ m[939] ^ m[941] ^ m[943] ^ m[945] ^ m[947] ^ m[949] ^ m[951] ^ m[953] ^ m[955] ^ m[957] ^ m[959] ^ m[960] ^ m[962] ^ m[964] ^ m[966] ^ m[968] ^ m[970] ^ m[972] ^ m[974] ^ m[976] ^ m[978] ^ m[980] ^ m[982] ^ m[984] ^ m[986] ^ m[988] ^ m[991] ^ m[993] ^ m[995] ^ m[997] ^ m[999] ^ m[1001] ^ m[1003] ^ m[1005] ^ m[1007] ^ m[1009] ^ m[1011] ^ m[1013] ^ m[1015] ^ m[1017] ^ m[1019] ^ m[1021] ^ m[1023] ^ m[1025] ^ m[1027] ^ m[1029] ^ m[1030] ^ m[1032] ^ m[1034] ^ m[1036] ^ m[1038] ^ m[1040] ^ m[1042] ^ m[1044] ^ m[1046] ^ m[1048] ^ m[1050] ^ m[1052] ^ m[1054] ^ m[1056] ^ m[1058] ^ m[1060] ^ m[1062] ^ m[1064] ^ m[1066] ^ m[1068] ^ m[1071] ^ m[1073] ^ m[1075] ^ m[1077] ^ m[1079] ^ m[1081] ^ m[1083] ^ m[1085] ^ m[1087] ^ m[1089] ^ m[1091] ^ m[1093] ^ m[1095] ^ m[1097] ^ m[1099] ^ m[1100] ^ m[1103] ^ m[1105] ^ m[1107] ^ m[1109] ^ m[1111] ^ m[1113] ^ m[1114] ^ m[1116] ^ m[1118] ^ m[1120] ^ m[1122] ^ m[1124] ^ m[1127] ^ m[1129] ^ m[1131] ^ m[1133] ^ m[1135] ^ m[1137] ^ m[1139] ^ m[1141] ^ m[1143] ^ m[1145] ^ m[1147] ^ m[1149] ^ m[1151] ^ m[1153] ^ m[1155] ^ m[1156] ^ m[1158] ^ m[1160] ^ m[1162] ^ m[1164] ^ m[1166] ^ m[1169] ^ m[1171] ^ m[1173] ^ m[1175] ^ m[1177] ^ m[1179] ^ m[1181] ^ m[1183] ^ m[1185] ^ m[1187] ^ m[1189] ^ m[1191] ^ m[1193] ^ m[1195] ^ m[1197] ^ m[1198] ^ m[1200] ^ m[1202] ^ m[1204] ^ m[1206] ^ m[1208] ^ m[1210] ^ m[1212] ^ m[1214] ^ m[1216] ^ m[1218] ^ m[1220] ^ m[1222] ^ m[1224] ^ m[1226] ^ m[1229] ^ m[1231] ^ m[1233] ^ m[1235] ^ m[1237] ^ m[1239] ^ m[1241] ^ m[1243] ^ m[1245] ^ m[1247] ^ m[1249] ^ m[1251] ^ m[1253] ^ m[1255] ^ m[1257] ^ m[1259] ^ m[1261] ^ m[1263] ^ m[1265] ^ m[1267] ^ m[1268] ^ m[1270] ^ m[1272] ^ m[1274] ^ m[1276] ^ m[1278] ^ m[1281] ^ m[1283] ^ m[1285] ^ m[1287] ^ m[1289] ^ m[1291] ^ m[1293] ^ m[1295] ^ m[1297] ^ m[1299] ^ m[1301] ^ m[1303] ^ m[1305] ^ m[1307] ^ m[1309] ^ m[1310] ^ m[1312] ^ m[1314] ^ m[1316] ^ m[1318] ^ m[1320] ^ m[1322] ^ m[1324] ^ m[1326] ^ m[1328] ^ m[1330] ^ m[1332] ^ m[1334] ^ m[1336] ^ m[1338] ^ m[1341] ^ m[1343] ^ m[1345] ^ m[1347] ^ m[1349] ^ m[1351] ^ m[1353] ^ m[1355] ^ m[1357] ^ m[1359] ^ m[1361] ^ m[1363] ^ m[1365] ^ m[1367] ^ m[1369] ^ m[1371] ^ m[1373] ^ m[1375] ^ m[1377] ^ m[1379] ^ m[1380] ^ m[1382] ^ m[1384] ^ m[1386] ^ m[1388] ^ m[1390] ^ m[1392] ^ m[1394] ^ m[1396] ^ m[1398] ^ m[1400] ^ m[1402] ^ m[1404] ^ m[1406] ^ m[1408] ^ m[1411] ^ m[1413] ^ m[1415] ^ m[1417] ^ m[1419] ^ m[1421] ^ m[1423] ^ m[1425] ^ m[1427] ^ m[1429] ^ m[1431] ^ m[1433] ^ m[1435] ^ m[1437] ^ m[1439] ^ m[1441] ^ m[1443] ^ m[1445] ^ m[1447] ^ m[1449] ^ m[1450] ^ m[1452] ^ m[1454] ^ m[1456] ^ m[1458] ^ m[1460] ^ m[1462] ^ m[1464] ^ m[1466] ^ m[1468] ^ m[1470] ^ m[1472] ^ m[1474] ^ m[1476] ^ m[1478] ^ m[1480] ^ m[1482] ^ m[1484] ^ m[1486] ^ m[1488] ^ m[1491] ^ m[1493] ^ m[1495] ^ m[1497] ^ m[1499] ^ m[1501] ^ m[1503] ^ m[1505] ^ m[1507] ^ m[1509] ^ m[1511] ^ m[1513] ^ m[1515] ^ m[1517] ^ m[1519] ^ m[1520] ^ m[1522] ^ m[1524] ^ m[1526] ^ m[1528] ^ m[1530] ^ m[1533] ^ m[1535] ^ m[1537] ^ m[1539] ^ m[1541] ^ m[1543] ^ m[1545] ^ m[1547] ^ m[1549] ^ m[1551] ^ m[1553] ^ m[1555] ^ m[1557] ^ m[1559] ^ m[1561] ^ m[1562] ^ m[1564] ^ m[1566] ^ m[1568] ^ m[1570] ^ m[1572] ^ m[1574] ^ m[1576] ^ m[1578] ^ m[1580] ^ m[1582] ^ m[1584] ^ m[1586] ^ m[1588] ^ m[1590] ^ m[1593] ^ m[1595] ^ m[1597] ^ m[1599] ^ m[1601] ^ m[1603] ^ m[1605] ^ m[1607] ^ m[1609] ^ m[1611] ^ m[1613] ^ m[1615] ^ m[1617] ^ m[1619] ^ m[1621] ^ m[1623] ^ m[1625] ^ m[1627] ^ m[1629] ^ m[1631] ^ m[1632] ^ m[1634] ^ m[1636] ^ m[1638] ^ m[1640] ^ m[1642] ^ m[1644] ^ m[1646] ^ m[1648] ^ m[1650] ^ m[1652] ^ m[1654] ^ m[1656] ^ m[1658] ^ m[1660] ^ m[1663] ^ m[1665] ^ m[1667] ^ m[1669] ^ m[1671] ^ m[1673] ^ m[1675] ^ m[1677] ^ m[1679] ^ m[1681] ^ m[1683] ^ m[1685] ^ m[1687] ^ m[1689] ^ m[1691] ^ m[1693] ^ m[1695] ^ m[1697] ^ m[1699] ^ m[1701] ^ m[1702] ^ m[1704] ^ m[1706] ^ m[1708] ^ m[1710] ^ m[1712] ^ m[1714] ^ m[1716] ^ m[1718] ^ m[1720] ^ m[1722] ^ m[1724] ^ m[1726] ^ m[1728] ^ m[1730] ^ m[1732] ^ m[1734] ^ m[1736] ^ m[1738] ^ m[1740] ^ m[1743] ^ m[1745] ^ m[1747] ^ m[1749] ^ m[1751] ^ m[1753] ^ m[1755] ^ m[1757] ^ m[1759] ^ m[1761] ^ m[1763] ^ m[1765] ^ m[1767] ^ m[1769] ^ m[1771] ^ m[1772] ^ m[1774] ^ m[1776] ^ m[1778] ^ m[1780] ^ m[1782] ^ m[1784] ^ m[1786] ^ m[1788] ^ m[1790] ^ m[1792] ^ m[1794] ^ m[1796] ^ m[1798] ^ m[1800] ^ m[1803] ^ m[1805] ^ m[1807] ^ m[1809] ^ m[1811] ^ m[1813] ^ m[1815] ^ m[1817] ^ m[1819] ^ m[1821] ^ m[1823] ^ m[1825] ^ m[1827] ^ m[1829] ^ m[1831] ^ m[1833] ^ m[1835] ^ m[1837] ^ m[1839] ^ m[1841] ^ m[1842] ^ m[1844] ^ m[1846] ^ m[1848] ^ m[1850] ^ m[1852] ^ m[1854] ^ m[1856] ^ m[1858] ^ m[1860] ^ m[1862] ^ m[1864] ^ m[1866] ^ m[1868] ^ m[1870] ^ m[1872] ^ m[1874] ^ m[1876] ^ m[1878] ^ m[1880] ^ m[1883] ^ m[1885] ^ m[1887] ^ m[1889] ^ m[1891] ^ m[1893] ^ m[1895] ^ m[1897] ^ m[1899] ^ m[1901] ^ m[1903] ^ m[1905] ^ m[1907] ^ m[1909] ^ m[1911] ^ m[1912] ^ m[1914] ^ m[1916] ^ m[1918] ^ m[1920] ^ m[1922] ^ m[1924] ^ m[1926] ^ m[1928] ^ m[1930] ^ m[1932] ^ m[1934] ^ m[1936] ^ m[1938] ^ m[1940] ^ m[1942] ^ m[1944] ^ m[1946] ^ m[1948] ^ m[1950] ^ m[1953] ^ m[1955] ^ m[1957] ^ m[1959] ^ m[1961] ^ m[1963] ^ m[1965] ^ m[1967] ^ m[1969] ^ m[1971] ^ m[1973] ^ m[1975] ^ m[1977] ^ m[1979] ^ m[1981] ^ m[1982] ^ m[1984] ^ m[1986] ^ m[1988] ^ m[1990] ^ m[1992] ^ m[1994] ^ m[1996] ^ m[1998] ^ m[2000] ^ m[2002] ^ m[2004] ^ m[2006] ^ m[2008] ^ m[2010] ^ m[2013] ^ m[2015] ^ m[2017] ^ m[2019] ^ m[2021] ^ m[2023] ^ m[2024] ^ m[2025] ^ m[2026] ^ m[2027] ^ m[2028] ^ m[2029] ^ m[2031] ^ m[2032] ^ m[2033] ^ m[2034] ^ m[2035];
    assign parity[7] = m[1] ^ m[3] ^ m[4] ^ m[7] ^ m[9] ^ m[11] ^ m[13] ^ m[15] ^ m[17] ^ m[19] ^ m[21] ^ m[22] ^ m[25] ^ m[27] ^ m[29] ^ m[31] ^ m[33] ^ m[35] ^ m[37] ^ m[38] ^ m[41] ^ m[43] ^ m[45] ^ m[47] ^ m[49] ^ m[51] ^ m[53] ^ m[54] ^ m[56] ^ m[58] ^ m[60] ^ m[62] ^ m[64] ^ m[66] ^ m[69] ^ m[71] ^ m[73] ^ m[75] ^ m[77] ^ m[79] ^ m[81] ^ m[83] ^ m[85] ^ m[87] ^ m[89] ^ m[91] ^ m[93] ^ m[95] ^ m[97] ^ m[99] ^ m[101] ^ m[103] ^ m[105] ^ m[107] ^ m[109] ^ m[111] ^ m[112] ^ m[115] ^ m[117] ^ m[119] ^ m[121] ^ m[123] ^ m[125] ^ m[127] ^ m[128] ^ m[131] ^ m[133] ^ m[135] ^ m[137] ^ m[139] ^ m[141] ^ m[143] ^ m[144] ^ m[146] ^ m[148] ^ m[150] ^ m[152] ^ m[154] ^ m[156] ^ m[159] ^ m[161] ^ m[163] ^ m[165] ^ m[167] ^ m[169] ^ m[171] ^ m[173] ^ m[175] ^ m[177] ^ m[179] ^ m[181] ^ m[183] ^ m[185] ^ m[187] ^ m[189] ^ m[191] ^ m[193] ^ m[195] ^ m[197] ^ m[199] ^ m[200] ^ m[203] ^ m[205] ^ m[207] ^ m[209] ^ m[211] ^ m[213] ^ m[215] ^ m[216] ^ m[218] ^ m[220] ^ m[222] ^ m[224] ^ m[226] ^ m[228] ^ m[231] ^ m[233] ^ m[235] ^ m[237] ^ m[239] ^ m[241] ^ m[243] ^ m[245] ^ m[247] ^ m[249] ^ m[251] ^ m[253] ^ m[255] ^ m[257] ^ m[259] ^ m[261] ^ m[263] ^ m[265] ^ m[267] ^ m[269] ^ m[271] ^ m[272] ^ m[274] ^ m[276] ^ m[278] ^ m[280] ^ m[282] ^ m[284] ^ m[287] ^ m[289] ^ m[291] ^ m[293] ^ m[295] ^ m[297] ^ m[299] ^ m[301] ^ m[303] ^ m[305] ^ m[307] ^ m[309] ^ m[311] ^ m[313] ^ m[315] ^ m[317] ^ m[319] ^ m[321] ^ m[323] ^ m[325] ^ m[327] ^ m[328] ^ m[330] ^ m[332] ^ m[334] ^ m[336] ^ m[338] ^ m[340] ^ m[342] ^ m[344] ^ m[346] ^ m[348] ^ m[350] ^ m[352] ^ m[354] ^ m[356] ^ m[358] ^ m[360] ^ m[362] ^ m[364] ^ m[366] ^ m[368] ^ m[371] ^ m[373] ^ m[375] ^ m[377] ^ m[379] ^ m[381] ^ m[383] ^ m[385] ^ m[387] ^ m[389] ^ m[391] ^ m[393] ^ m[395] ^ m[397] ^ m[399] ^ m[401] ^ m[403] ^ m[405] ^ m[407] ^ m[409] ^ m[411] ^ m[413] ^ m[415] ^ m[417] ^ m[419] ^ m[421] ^ m[423] ^ m[425] ^ m[427] ^ m[429] ^ m[431] ^ m[433] ^ m[435] ^ m[437] ^ m[439] ^ m[440] ^ m[443] ^ m[445] ^ m[447] ^ m[449] ^ m[451] ^ m[453] ^ m[455] ^ m[456] ^ m[458] ^ m[460] ^ m[462] ^ m[464] ^ m[466] ^ m[468] ^ m[471] ^ m[473] ^ m[475] ^ m[477] ^ m[479] ^ m[481] ^ m[483] ^ m[485] ^ m[487] ^ m[489] ^ m[491] ^ m[493] ^ m[495] ^ m[497] ^ m[499] ^ m[501] ^ m[503] ^ m[505] ^ m[507] ^ m[509] ^ m[511] ^ m[512] ^ m[514] ^ m[516] ^ m[518] ^ m[520] ^ m[522] ^ m[524] ^ m[527] ^ m[529] ^ m[531] ^ m[533] ^ m[535] ^ m[537] ^ m[539] ^ m[541] ^ m[543] ^ m[545] ^ m[547] ^ m[549] ^ m[551] ^ m[553] ^ m[555] ^ m[557] ^ m[559] ^ m[561] ^ m[563] ^ m[565] ^ m[567] ^ m[568] ^ m[570] ^ m[572] ^ m[574] ^ m[576] ^ m[578] ^ m[580] ^ m[582] ^ m[584] ^ m[586] ^ m[588] ^ m[590] ^ m[592] ^ m[594] ^ m[596] ^ m[598] ^ m[600] ^ m[602] ^ m[604] ^ m[606] ^ m[608] ^ m[611] ^ m[613] ^ m[615] ^ m[617] ^ m[619] ^ m[621] ^ m[623] ^ m[625] ^ m[627] ^ m[629] ^ m[631] ^ m[633] ^ m[635] ^ m[637] ^ m[639] ^ m[641] ^ m[643] ^ m[645] ^ m[647] ^ m[649] ^ m[651] ^ m[653] ^ m[655] ^ m[657] ^ m[659] ^ m[661] ^ m[663] ^ m[665] ^ m[667] ^ m[669] ^ m[671] ^ m[673] ^ m[675] ^ m[677] ^ m[679] ^ m[680] ^ m[682] ^ m[684] ^ m[686] ^ m[688] ^ m[690] ^ m[692] ^ m[695] ^ m[697] ^ m[699] ^ m[701] ^ m[703] ^ m[705] ^ m[707] ^ m[709] ^ m[711] ^ m[713] ^ m[715] ^ m[717] ^ m[719] ^ m[721] ^ m[723] ^ m[725] ^ m[727] ^ m[729] ^ m[731] ^ m[733] ^ m[735] ^ m[736] ^ m[738] ^ m[740] ^ m[742] ^ m[744] ^ m[746] ^ m[748] ^ m[750] ^ m[752] ^ m[754] ^ m[756] ^ m[758] ^ m[760] ^ m[762] ^ m[764] ^ m[766] ^ m[768] ^ m[770] ^ m[772] ^ m[774] ^ m[776] ^ m[779] ^ m[781] ^ m[783] ^ m[785] ^ m[787] ^ m[789] ^ m[791] ^ m[793] ^ m[795] ^ m[797] ^ m[799] ^ m[801] ^ m[803] ^ m[805] ^ m[807] ^ m[809] ^ m[811] ^ m[813] ^ m[815] ^ m[817] ^ m[819] ^ m[821] ^ m[823] ^ m[825] ^ m[827] ^ m[829] ^ m[831] ^ m[833] ^ m[835] ^ m[837] ^ m[839] ^ m[841] ^ m[843] ^ m[845] ^ m[847] ^ m[848] ^ m[850] ^ m[852] ^ m[854] ^ m[856] ^ m[858] ^ m[860] ^ m[862] ^ m[864] ^ m[866] ^ m[868] ^ m[870] ^ m[872] ^ m[874] ^ m[876] ^ m[878] ^ m[880] ^ m[882] ^ m[884] ^ m[886] ^ m[888] ^ m[891] ^ m[893] ^ m[895] ^ m[897] ^ m[899] ^ m[901] ^ m[903] ^ m[905] ^ m[907] ^ m[909] ^ m[911] ^ m[913] ^ m[915] ^ m[917] ^ m[919] ^ m[921] ^ m[923] ^ m[925] ^ m[927] ^ m[929] ^ m[931] ^ m[933] ^ m[935] ^ m[937] ^ m[939] ^ m[941] ^ m[943] ^ m[945] ^ m[947] ^ m[949] ^ m[951] ^ m[953] ^ m[955] ^ m[957] ^ m[959] ^ m[960] ^ m[962] ^ m[964] ^ m[966] ^ m[968] ^ m[970] ^ m[972] ^ m[974] ^ m[976] ^ m[978] ^ m[980] ^ m[982] ^ m[984] ^ m[986] ^ m[988] ^ m[990] ^ m[992] ^ m[994] ^ m[996] ^ m[998] ^ m[1000] ^ m[1002] ^ m[1004] ^ m[1006] ^ m[1008] ^ m[1010] ^ m[1012] ^ m[1014] ^ m[1016] ^ m[1018] ^ m[1020] ^ m[1022] ^ m[1024] ^ m[1026] ^ m[1028] ^ m[1031] ^ m[1033] ^ m[1035] ^ m[1037] ^ m[1039] ^ m[1041] ^ m[1043] ^ m[1045] ^ m[1047] ^ m[1049] ^ m[1051] ^ m[1053] ^ m[1055] ^ m[1057] ^ m[1059] ^ m[1061] ^ m[1063] ^ m[1065] ^ m[1067] ^ m[1069] ^ m[1071] ^ m[1073] ^ m[1075] ^ m[1077] ^ m[1079] ^ m[1081] ^ m[1083] ^ m[1085] ^ m[1087] ^ m[1089] ^ m[1091] ^ m[1093] ^ m[1095] ^ m[1097] ^ m[1099] ^ m[1100] ^ m[1102] ^ m[1104] ^ m[1106] ^ m[1108] ^ m[1110] ^ m[1112] ^ m[1115] ^ m[1117] ^ m[1119] ^ m[1121] ^ m[1123] ^ m[1125] ^ m[1127] ^ m[1129] ^ m[1131] ^ m[1133] ^ m[1135] ^ m[1137] ^ m[1139] ^ m[1141] ^ m[1143] ^ m[1145] ^ m[1147] ^ m[1149] ^ m[1151] ^ m[1153] ^ m[1155] ^ m[1156] ^ m[1158] ^ m[1160] ^ m[1162] ^ m[1164] ^ m[1166] ^ m[1168] ^ m[1170] ^ m[1172] ^ m[1174] ^ m[1176] ^ m[1178] ^ m[1180] ^ m[1182] ^ m[1184] ^ m[1186] ^ m[1188] ^ m[1190] ^ m[1192] ^ m[1194] ^ m[1196] ^ m[1199] ^ m[1201] ^ m[1203] ^ m[1205] ^ m[1207] ^ m[1209] ^ m[1211] ^ m[1213] ^ m[1215] ^ m[1217] ^ m[1219] ^ m[1221] ^ m[1223] ^ m[1225] ^ m[1227] ^ m[1229] ^ m[1231] ^ m[1233] ^ m[1235] ^ m[1237] ^ m[1239] ^ m[1241] ^ m[1243] ^ m[1245] ^ m[1247] ^ m[1249] ^ m[1251] ^ m[1253] ^ m[1255] ^ m[1257] ^ m[1259] ^ m[1261] ^ m[1263] ^ m[1265] ^ m[1267] ^ m[1268] ^ m[1270] ^ m[1272] ^ m[1274] ^ m[1276] ^ m[1278] ^ m[1280] ^ m[1282] ^ m[1284] ^ m[1286] ^ m[1288] ^ m[1290] ^ m[1292] ^ m[1294] ^ m[1296] ^ m[1298] ^ m[1300] ^ m[1302] ^ m[1304] ^ m[1306] ^ m[1308] ^ m[1311] ^ m[1313] ^ m[1315] ^ m[1317] ^ m[1319] ^ m[1321] ^ m[1323] ^ m[1325] ^ m[1327] ^ m[1329] ^ m[1331] ^ m[1333] ^ m[1335] ^ m[1337] ^ m[1339] ^ m[1341] ^ m[1343] ^ m[1345] ^ m[1347] ^ m[1349] ^ m[1351] ^ m[1353] ^ m[1355] ^ m[1357] ^ m[1359] ^ m[1361] ^ m[1363] ^ m[1365] ^ m[1367] ^ m[1369] ^ m[1371] ^ m[1373] ^ m[1375] ^ m[1377] ^ m[1379] ^ m[1380] ^ m[1382] ^ m[1384] ^ m[1386] ^ m[1388] ^ m[1390] ^ m[1392] ^ m[1394] ^ m[1396] ^ m[1398] ^ m[1400] ^ m[1402] ^ m[1404] ^ m[1406] ^ m[1408] ^ m[1410] ^ m[1412] ^ m[1414] ^ m[1416] ^ m[1418] ^ m[1420] ^ m[1422] ^ m[1424] ^ m[1426] ^ m[1428] ^ m[1430] ^ m[1432] ^ m[1434] ^ m[1436] ^ m[1438] ^ m[1440] ^ m[1442] ^ m[1444] ^ m[1446] ^ m[1448] ^ m[1451] ^ m[1453] ^ m[1455] ^ m[1457] ^ m[1459] ^ m[1461] ^ m[1463] ^ m[1465] ^ m[1467] ^ m[1469] ^ m[1471] ^ m[1473] ^ m[1475] ^ m[1477] ^ m[1479] ^ m[1481] ^ m[1483] ^ m[1485] ^ m[1487] ^ m[1489] ^ m[1491] ^ m[1493] ^ m[1495] ^ m[1497] ^ m[1499] ^ m[1501] ^ m[1503] ^ m[1505] ^ m[1507] ^ m[1509] ^ m[1511] ^ m[1513] ^ m[1515] ^ m[1517] ^ m[1519] ^ m[1520] ^ m[1522] ^ m[1524] ^ m[1526] ^ m[1528] ^ m[1530] ^ m[1532] ^ m[1534] ^ m[1536] ^ m[1538] ^ m[1540] ^ m[1542] ^ m[1544] ^ m[1546] ^ m[1548] ^ m[1550] ^ m[1552] ^ m[1554] ^ m[1556] ^ m[1558] ^ m[1560] ^ m[1563] ^ m[1565] ^ m[1567] ^ m[1569] ^ m[1571] ^ m[1573] ^ m[1575] ^ m[1577] ^ m[1579] ^ m[1581] ^ m[1583] ^ m[1585] ^ m[1587] ^ m[1589] ^ m[1591] ^ m[1593] ^ m[1595] ^ m[1597] ^ m[1599] ^ m[1601] ^ m[1603] ^ m[1605] ^ m[1607] ^ m[1609] ^ m[1611] ^ m[1613] ^ m[1615] ^ m[1617] ^ m[1619] ^ m[1621] ^ m[1623] ^ m[1625] ^ m[1627] ^ m[1629] ^ m[1631] ^ m[1632] ^ m[1634] ^ m[1636] ^ m[1638] ^ m[1640] ^ m[1642] ^ m[1644] ^ m[1646] ^ m[1648] ^ m[1650] ^ m[1652] ^ m[1654] ^ m[1656] ^ m[1658] ^ m[1660] ^ m[1662] ^ m[1664] ^ m[1666] ^ m[1668] ^ m[1670] ^ m[1672] ^ m[1674] ^ m[1676] ^ m[1678] ^ m[1680] ^ m[1682] ^ m[1684] ^ m[1686] ^ m[1688] ^ m[1690] ^ m[1692] ^ m[1694] ^ m[1696] ^ m[1698] ^ m[1700] ^ m[1703] ^ m[1705] ^ m[1707] ^ m[1709] ^ m[1711] ^ m[1713] ^ m[1715] ^ m[1717] ^ m[1719] ^ m[1721] ^ m[1723] ^ m[1725] ^ m[1727] ^ m[1729] ^ m[1731] ^ m[1733] ^ m[1735] ^ m[1737] ^ m[1739] ^ m[1741] ^ m[1743] ^ m[1745] ^ m[1747] ^ m[1749] ^ m[1751] ^ m[1753] ^ m[1755] ^ m[1757] ^ m[1759] ^ m[1761] ^ m[1763] ^ m[1765] ^ m[1767] ^ m[1769] ^ m[1771] ^ m[1772] ^ m[1774] ^ m[1776] ^ m[1778] ^ m[1780] ^ m[1782] ^ m[1784] ^ m[1786] ^ m[1788] ^ m[1790] ^ m[1792] ^ m[1794] ^ m[1796] ^ m[1798] ^ m[1800] ^ m[1802] ^ m[1804] ^ m[1806] ^ m[1808] ^ m[1810] ^ m[1812] ^ m[1814] ^ m[1816] ^ m[1818] ^ m[1820] ^ m[1822] ^ m[1824] ^ m[1826] ^ m[1828] ^ m[1830] ^ m[1832] ^ m[1834] ^ m[1836] ^ m[1838] ^ m[1840] ^ m[1843] ^ m[1845] ^ m[1847] ^ m[1849] ^ m[1851] ^ m[1853] ^ m[1855] ^ m[1857] ^ m[1859] ^ m[1861] ^ m[1863] ^ m[1865] ^ m[1867] ^ m[1869] ^ m[1871] ^ m[1873] ^ m[1875] ^ m[1877] ^ m[1879] ^ m[1881] ^ m[1883] ^ m[1885] ^ m[1887] ^ m[1889] ^ m[1891] ^ m[1893] ^ m[1895] ^ m[1897] ^ m[1899] ^ m[1901] ^ m[1903] ^ m[1905] ^ m[1907] ^ m[1909] ^ m[1911] ^ m[1912] ^ m[1914] ^ m[1916] ^ m[1918] ^ m[1920] ^ m[1922] ^ m[1924] ^ m[1926] ^ m[1928] ^ m[1930] ^ m[1932] ^ m[1934] ^ m[1936] ^ m[1938] ^ m[1940] ^ m[1942] ^ m[1944] ^ m[1946] ^ m[1948] ^ m[1950] ^ m[1952] ^ m[1954] ^ m[1956] ^ m[1958] ^ m[1960] ^ m[1962] ^ m[1964] ^ m[1966] ^ m[1968] ^ m[1970] ^ m[1972] ^ m[1974] ^ m[1976] ^ m[1978] ^ m[1980] ^ m[1983] ^ m[1985] ^ m[1987] ^ m[1989] ^ m[1991] ^ m[1993] ^ m[1995] ^ m[1997] ^ m[1999] ^ m[2001] ^ m[2003] ^ m[2005] ^ m[2007] ^ m[2009] ^ m[2011] ^ m[2013] ^ m[2015] ^ m[2017] ^ m[2019] ^ m[2021] ^ m[2023] ^ m[2024] ^ m[2025] ^ m[2026] ^ m[2027] ^ m[2028] ^ m[2029] ^ m[2030] ^ m[2032] ^ m[2033] ^ m[2034] ^ m[2035];
    assign parity[8] = m[1] ^ m[2] ^ m[5] ^ m[7] ^ m[9] ^ m[11] ^ m[13] ^ m[15] ^ m[17] ^ m[19] ^ m[20] ^ m[23] ^ m[25] ^ m[27] ^ m[29] ^ m[31] ^ m[33] ^ m[35] ^ m[37] ^ m[38] ^ m[40] ^ m[42] ^ m[44] ^ m[46] ^ m[48] ^ m[50] ^ m[52] ^ m[55] ^ m[57] ^ m[59] ^ m[61] ^ m[63] ^ m[65] ^ m[67] ^ m[69] ^ m[71] ^ m[73] ^ m[75] ^ m[77] ^ m[79] ^ m[81] ^ m[83] ^ m[85] ^ m[87] ^ m[89] ^ m[91] ^ m[93] ^ m[95] ^ m[97] ^ m[99] ^ m[101] ^ m[103] ^ m[105] ^ m[107] ^ m[109] ^ m[110] ^ m[113] ^ m[115] ^ m[117] ^ m[119] ^ m[121] ^ m[123] ^ m[125] ^ m[127] ^ m[128] ^ m[130] ^ m[132] ^ m[134] ^ m[136] ^ m[138] ^ m[140] ^ m[142] ^ m[145] ^ m[147] ^ m[149] ^ m[151] ^ m[153] ^ m[155] ^ m[157] ^ m[159] ^ m[161] ^ m[163] ^ m[165] ^ m[167] ^ m[169] ^ m[171] ^ m[173] ^ m[175] ^ m[177] ^ m[179] ^ m[181] ^ m[183] ^ m[185] ^ m[187] ^ m[189] ^ m[191] ^ m[193] ^ m[195] ^ m[197] ^ m[199] ^ m[200] ^ m[202] ^ m[204] ^ m[206] ^ m[208] ^ m[210] ^ m[212] ^ m[214] ^ m[217] ^ m[219] ^ m[221] ^ m[223] ^ m[225] ^ m[227] ^ m[229] ^ m[231] ^ m[233] ^ m[235] ^ m[237] ^ m[239] ^ m[241] ^ m[243] ^ m[245] ^ m[247] ^ m[249] ^ m[251] ^ m[253] ^ m[255] ^ m[257] ^ m[259] ^ m[261] ^ m[263] ^ m[265] ^ m[267] ^ m[269] ^ m[271] ^ m[272] ^ m[274] ^ m[276] ^ m[278] ^ m[280] ^ m[282] ^ m[284] ^ m[286] ^ m[288] ^ m[290] ^ m[292] ^ m[294] ^ m[296] ^ m[298] ^ m[300] ^ m[302] ^ m[304] ^ m[306] ^ m[308] ^ m[310] ^ m[312] ^ m[314] ^ m[316] ^ m[318] ^ m[320] ^ m[322] ^ m[324] ^ m[326] ^ m[329] ^ m[331] ^ m[333] ^ m[335] ^ m[337] ^ m[339] ^ m[341] ^ m[343] ^ m[345] ^ m[347] ^ m[349] ^ m[351] ^ m[353] ^ m[355] ^ m[357] ^ m[359] ^ m[361] ^ m[363] ^ m[365] ^ m[367] ^ m[369] ^ m[371] ^ m[373] ^ m[375] ^ m[377] ^ m[379] ^ m[381] ^ m[383] ^ m[385] ^ m[387] ^ m[389] ^ m[391] ^ m[393] ^ m[395] ^ m[397] ^ m[399] ^ m[401] ^ m[403] ^ m[405] ^ m[407] ^ m[409] ^ m[411] ^ m[413] ^ m[415] ^ m[417] ^ m[419] ^ m[421] ^ m[423] ^ m[425] ^ m[427] ^ m[429] ^ m[431] ^ m[433] ^ m[435] ^ m[437] ^ m[439] ^ m[440] ^ m[442] ^ m[444] ^ m[446] ^ m[448] ^ m[450] ^ m[452] ^ m[454] ^ m[457] ^ m[459] ^ m[461] ^ m[463] ^ m[465] ^ m[467] ^ m[469] ^ m[471] ^ m[473] ^ m[475] ^ m[477] ^ m[479] ^ m[481] ^ m[483] ^ m[485] ^ m[487] ^ m[489] ^ m[491] ^ m[493] ^ m[495] ^ m[497] ^ m[499] ^ m[501] ^ m[503] ^ m[505] ^ m[507] ^ m[509] ^ m[511] ^ m[512] ^ m[514] ^ m[516] ^ m[518] ^ m[520] ^ m[522] ^ m[524] ^ m[526] ^ m[528] ^ m[530] ^ m[532] ^ m[534] ^ m[536] ^ m[538] ^ m[540] ^ m[542] ^ m[544] ^ m[546] ^ m[548] ^ m[550] ^ m[552] ^ m[554] ^ m[556] ^ m[558] ^ m[560] ^ m[562] ^ m[564] ^ m[566] ^ m[569] ^ m[571] ^ m[573] ^ m[575] ^ m[577] ^ m[579] ^ m[581] ^ m[583] ^ m[585] ^ m[587] ^ m[589] ^ m[591] ^ m[593] ^ m[595] ^ m[597] ^ m[599] ^ m[601] ^ m[603] ^ m[605] ^ m[607] ^ m[609] ^ m[611] ^ m[613] ^ m[615] ^ m[617] ^ m[619] ^ m[621] ^ m[623] ^ m[625] ^ m[627] ^ m[629] ^ m[631] ^ m[633] ^ m[635] ^ m[637] ^ m[639] ^ m[641] ^ m[643] ^ m[645] ^ m[647] ^ m[649] ^ m[651] ^ m[653] ^ m[655] ^ m[657] ^ m[659] ^ m[661] ^ m[663] ^ m[665] ^ m[667] ^ m[669] ^ m[671] ^ m[673] ^ m[675] ^ m[677] ^ m[679] ^ m[680] ^ m[682] ^ m[684] ^ m[686] ^ m[688] ^ m[690] ^ m[692] ^ m[694] ^ m[696] ^ m[698] ^ m[700] ^ m[702] ^ m[704] ^ m[706] ^ m[708] ^ m[710] ^ m[712] ^ m[714] ^ m[716] ^ m[718] ^ m[720] ^ m[722] ^ m[724] ^ m[726] ^ m[728] ^ m[730] ^ m[732] ^ m[734] ^ m[737] ^ m[739] ^ m[741] ^ m[743] ^ m[745] ^ m[747] ^ m[749] ^ m[751] ^ m[753] ^ m[755] ^ m[757] ^ m[759] ^ m[761] ^ m[763] ^ m[765] ^ m[767] ^ m[769] ^ m[771] ^ m[773] ^ m[775] ^ m[777] ^ m[779] ^ m[781] ^ m[783] ^ m[785] ^ m[787] ^ m[789] ^ m[791] ^ m[793] ^ m[795] ^ m[797] ^ m[799] ^ m[801] ^ m[803] ^ m[805] ^ m[807] ^ m[809] ^ m[811] ^ m[813] ^ m[815] ^ m[817] ^ m[819] ^ m[821] ^ m[823] ^ m[825] ^ m[827] ^ m[829] ^ m[831] ^ m[833] ^ m[835] ^ m[837] ^ m[839] ^ m[841] ^ m[843] ^ m[845] ^ m[847] ^ m[848] ^ m[850] ^ m[852] ^ m[854] ^ m[856] ^ m[858] ^ m[860] ^ m[862] ^ m[864] ^ m[866] ^ m[868] ^ m[870] ^ m[872] ^ m[874] ^ m[876] ^ m[878] ^ m[880] ^ m[882] ^ m[884] ^ m[886] ^ m[888] ^ m[890] ^ m[892] ^ m[894] ^ m[896] ^ m[898] ^ m[900] ^ m[902] ^ m[904] ^ m[906] ^ m[908] ^ m[910] ^ m[912] ^ m[914] ^ m[916] ^ m[918] ^ m[920] ^ m[922] ^ m[924] ^ m[926] ^ m[928] ^ m[930] ^ m[932] ^ m[934] ^ m[936] ^ m[938] ^ m[940] ^ m[942] ^ m[944] ^ m[946] ^ m[948] ^ m[950] ^ m[952] ^ m[954] ^ m[956] ^ m[958] ^ m[961] ^ m[963] ^ m[965] ^ m[967] ^ m[969] ^ m[971] ^ m[973] ^ m[975] ^ m[977] ^ m[979] ^ m[981] ^ m[983] ^ m[985] ^ m[987] ^ m[989] ^ m[991] ^ m[993] ^ m[995] ^ m[997] ^ m[999] ^ m[1001] ^ m[1003] ^ m[1005] ^ m[1007] ^ m[1009] ^ m[1011] ^ m[1013] ^ m[1015] ^ m[1017] ^ m[1019] ^ m[1021] ^ m[1023] ^ m[1025] ^ m[1027] ^ m[1029] ^ m[1031] ^ m[1033] ^ m[1035] ^ m[1037] ^ m[1039] ^ m[1041] ^ m[1043] ^ m[1045] ^ m[1047] ^ m[1049] ^ m[1051] ^ m[1053] ^ m[1055] ^ m[1057] ^ m[1059] ^ m[1061] ^ m[1063] ^ m[1065] ^ m[1067] ^ m[1069] ^ m[1071] ^ m[1073] ^ m[1075] ^ m[1077] ^ m[1079] ^ m[1081] ^ m[1083] ^ m[1085] ^ m[1087] ^ m[1089] ^ m[1091] ^ m[1093] ^ m[1095] ^ m[1097] ^ m[1099] ^ m[1100] ^ m[1102] ^ m[1104] ^ m[1106] ^ m[1108] ^ m[1110] ^ m[1112] ^ m[1114] ^ m[1116] ^ m[1118] ^ m[1120] ^ m[1122] ^ m[1124] ^ m[1126] ^ m[1128] ^ m[1130] ^ m[1132] ^ m[1134] ^ m[1136] ^ m[1138] ^ m[1140] ^ m[1142] ^ m[1144] ^ m[1146] ^ m[1148] ^ m[1150] ^ m[1152] ^ m[1154] ^ m[1157] ^ m[1159] ^ m[1161] ^ m[1163] ^ m[1165] ^ m[1167] ^ m[1169] ^ m[1171] ^ m[1173] ^ m[1175] ^ m[1177] ^ m[1179] ^ m[1181] ^ m[1183] ^ m[1185] ^ m[1187] ^ m[1189] ^ m[1191] ^ m[1193] ^ m[1195] ^ m[1197] ^ m[1199] ^ m[1201] ^ m[1203] ^ m[1205] ^ m[1207] ^ m[1209] ^ m[1211] ^ m[1213] ^ m[1215] ^ m[1217] ^ m[1219] ^ m[1221] ^ m[1223] ^ m[1225] ^ m[1227] ^ m[1229] ^ m[1231] ^ m[1233] ^ m[1235] ^ m[1237] ^ m[1239] ^ m[1241] ^ m[1243] ^ m[1245] ^ m[1247] ^ m[1249] ^ m[1251] ^ m[1253] ^ m[1255] ^ m[1257] ^ m[1259] ^ m[1261] ^ m[1263] ^ m[1265] ^ m[1267] ^ m[1268] ^ m[1270] ^ m[1272] ^ m[1274] ^ m[1276] ^ m[1278] ^ m[1280] ^ m[1282] ^ m[1284] ^ m[1286] ^ m[1288] ^ m[1290] ^ m[1292] ^ m[1294] ^ m[1296] ^ m[1298] ^ m[1300] ^ m[1302] ^ m[1304] ^ m[1306] ^ m[1308] ^ m[1310] ^ m[1312] ^ m[1314] ^ m[1316] ^ m[1318] ^ m[1320] ^ m[1322] ^ m[1324] ^ m[1326] ^ m[1328] ^ m[1330] ^ m[1332] ^ m[1334] ^ m[1336] ^ m[1338] ^ m[1340] ^ m[1342] ^ m[1344] ^ m[1346] ^ m[1348] ^ m[1350] ^ m[1352] ^ m[1354] ^ m[1356] ^ m[1358] ^ m[1360] ^ m[1362] ^ m[1364] ^ m[1366] ^ m[1368] ^ m[1370] ^ m[1372] ^ m[1374] ^ m[1376] ^ m[1378] ^ m[1381] ^ m[1383] ^ m[1385] ^ m[1387] ^ m[1389] ^ m[1391] ^ m[1393] ^ m[1395] ^ m[1397] ^ m[1399] ^ m[1401] ^ m[1403] ^ m[1405] ^ m[1407] ^ m[1409] ^ m[1411] ^ m[1413] ^ m[1415] ^ m[1417] ^ m[1419] ^ m[1421] ^ m[1423] ^ m[1425] ^ m[1427] ^ m[1429] ^ m[1431] ^ m[1433] ^ m[1435] ^ m[1437] ^ m[1439] ^ m[1441] ^ m[1443] ^ m[1445] ^ m[1447] ^ m[1449] ^ m[1451] ^ m[1453] ^ m[1455] ^ m[1457] ^ m[1459] ^ m[1461] ^ m[1463] ^ m[1465] ^ m[1467] ^ m[1469] ^ m[1471] ^ m[1473] ^ m[1475] ^ m[1477] ^ m[1479] ^ m[1481] ^ m[1483] ^ m[1485] ^ m[1487] ^ m[1489] ^ m[1491] ^ m[1493] ^ m[1495] ^ m[1497] ^ m[1499] ^ m[1501] ^ m[1503] ^ m[1505] ^ m[1507] ^ m[1509] ^ m[1511] ^ m[1513] ^ m[1515] ^ m[1517] ^ m[1519] ^ m[1520] ^ m[1522] ^ m[1524] ^ m[1526] ^ m[1528] ^ m[1530] ^ m[1532] ^ m[1534] ^ m[1536] ^ m[1538] ^ m[1540] ^ m[1542] ^ m[1544] ^ m[1546] ^ m[1548] ^ m[1550] ^ m[1552] ^ m[1554] ^ m[1556] ^ m[1558] ^ m[1560] ^ m[1562] ^ m[1564] ^ m[1566] ^ m[1568] ^ m[1570] ^ m[1572] ^ m[1574] ^ m[1576] ^ m[1578] ^ m[1580] ^ m[1582] ^ m[1584] ^ m[1586] ^ m[1588] ^ m[1590] ^ m[1592] ^ m[1594] ^ m[1596] ^ m[1598] ^ m[1600] ^ m[1602] ^ m[1604] ^ m[1606] ^ m[1608] ^ m[1610] ^ m[1612] ^ m[1614] ^ m[1616] ^ m[1618] ^ m[1620] ^ m[1622] ^ m[1624] ^ m[1626] ^ m[1628] ^ m[1630] ^ m[1633] ^ m[1635] ^ m[1637] ^ m[1639] ^ m[1641] ^ m[1643] ^ m[1645] ^ m[1647] ^ m[1649] ^ m[1651] ^ m[1653] ^ m[1655] ^ m[1657] ^ m[1659] ^ m[1661] ^ m[1663] ^ m[1665] ^ m[1667] ^ m[1669] ^ m[1671] ^ m[1673] ^ m[1675] ^ m[1677] ^ m[1679] ^ m[1681] ^ m[1683] ^ m[1685] ^ m[1687] ^ m[1689] ^ m[1691] ^ m[1693] ^ m[1695] ^ m[1697] ^ m[1699] ^ m[1701] ^ m[1703] ^ m[1705] ^ m[1707] ^ m[1709] ^ m[1711] ^ m[1713] ^ m[1715] ^ m[1717] ^ m[1719] ^ m[1721] ^ m[1723] ^ m[1725] ^ m[1727] ^ m[1729] ^ m[1731] ^ m[1733] ^ m[1735] ^ m[1737] ^ m[1739] ^ m[1741] ^ m[1743] ^ m[1745] ^ m[1747] ^ m[1749] ^ m[1751] ^ m[1753] ^ m[1755] ^ m[1757] ^ m[1759] ^ m[1761] ^ m[1763] ^ m[1765] ^ m[1767] ^ m[1769] ^ m[1771] ^ m[1772] ^ m[1774] ^ m[1776] ^ m[1778] ^ m[1780] ^ m[1782] ^ m[1784] ^ m[1786] ^ m[1788] ^ m[1790] ^ m[1792] ^ m[1794] ^ m[1796] ^ m[1798] ^ m[1800] ^ m[1802] ^ m[1804] ^ m[1806] ^ m[1808] ^ m[1810] ^ m[1812] ^ m[1814] ^ m[1816] ^ m[1818] ^ m[1820] ^ m[1822] ^ m[1824] ^ m[1826] ^ m[1828] ^ m[1830] ^ m[1832] ^ m[1834] ^ m[1836] ^ m[1838] ^ m[1840] ^ m[1842] ^ m[1844] ^ m[1846] ^ m[1848] ^ m[1850] ^ m[1852] ^ m[1854] ^ m[1856] ^ m[1858] ^ m[1860] ^ m[1862] ^ m[1864] ^ m[1866] ^ m[1868] ^ m[1870] ^ m[1872] ^ m[1874] ^ m[1876] ^ m[1878] ^ m[1880] ^ m[1882] ^ m[1884] ^ m[1886] ^ m[1888] ^ m[1890] ^ m[1892] ^ m[1894] ^ m[1896] ^ m[1898] ^ m[1900] ^ m[1902] ^ m[1904] ^ m[1906] ^ m[1908] ^ m[1910] ^ m[1913] ^ m[1915] ^ m[1917] ^ m[1919] ^ m[1921] ^ m[1923] ^ m[1925] ^ m[1927] ^ m[1929] ^ m[1931] ^ m[1933] ^ m[1935] ^ m[1937] ^ m[1939] ^ m[1941] ^ m[1943] ^ m[1945] ^ m[1947] ^ m[1949] ^ m[1951] ^ m[1953] ^ m[1955] ^ m[1957] ^ m[1959] ^ m[1961] ^ m[1963] ^ m[1965] ^ m[1967] ^ m[1969] ^ m[1971] ^ m[1973] ^ m[1975] ^ m[1977] ^ m[1979] ^ m[1981] ^ m[1983] ^ m[1985] ^ m[1987] ^ m[1989] ^ m[1991] ^ m[1993] ^ m[1995] ^ m[1997] ^ m[1999] ^ m[2001] ^ m[2003] ^ m[2005] ^ m[2007] ^ m[2009] ^ m[2011] ^ m[2013] ^ m[2015] ^ m[2017] ^ m[2019] ^ m[2021] ^ m[2023] ^ m[2024] ^ m[2025] ^ m[2026] ^ m[2027] ^ m[2028] ^ m[2029] ^ m[2030] ^ m[2031] ^ m[2033] ^ m[2034] ^ m[2035];
    assign parity[9] = m[0] ^ m[3] ^ m[5] ^ m[7] ^ m[9] ^ m[11] ^ m[13] ^ m[15] ^ m[17] ^ m[19] ^ m[20] ^ m[22] ^ m[24] ^ m[26] ^ m[28] ^ m[30] ^ m[32] ^ m[34] ^ m[36] ^ m[39] ^ m[41] ^ m[43] ^ m[45] ^ m[47] ^ m[49] ^ m[51] ^ m[53] ^ m[55] ^ m[57] ^ m[59] ^ m[61] ^ m[63] ^ m[65] ^ m[67] ^ m[69] ^ m[71] ^ m[73] ^ m[75] ^ m[77] ^ m[79] ^ m[81] ^ m[83] ^ m[85] ^ m[87] ^ m[89] ^ m[91] ^ m[93] ^ m[95] ^ m[97] ^ m[99] ^ m[101] ^ m[103] ^ m[105] ^ m[107] ^ m[109] ^ m[110] ^ m[112] ^ m[114] ^ m[116] ^ m[118] ^ m[120] ^ m[122] ^ m[124] ^ m[126] ^ m[129] ^ m[131] ^ m[133] ^ m[135] ^ m[137] ^ m[139] ^ m[141] ^ m[143] ^ m[145] ^ m[147] ^ m[149] ^ m[151] ^ m[153] ^ m[155] ^ m[157] ^ m[159] ^ m[161] ^ m[163] ^ m[165] ^ m[167] ^ m[169] ^ m[171] ^ m[173] ^ m[175] ^ m[177] ^ m[179] ^ m[181] ^ m[183] ^ m[185] ^ m[187] ^ m[189] ^ m[191] ^ m[193] ^ m[195] ^ m[197] ^ m[199] ^ m[200] ^ m[202] ^ m[204] ^ m[206] ^ m[208] ^ m[210] ^ m[212] ^ m[214] ^ m[216] ^ m[218] ^ m[220] ^ m[222] ^ m[224] ^ m[226] ^ m[228] ^ m[230] ^ m[232] ^ m[234] ^ m[236] ^ m[238] ^ m[240] ^ m[242] ^ m[244] ^ m[246] ^ m[248] ^ m[250] ^ m[252] ^ m[254] ^ m[256] ^ m[258] ^ m[260] ^ m[262] ^ m[264] ^ m[266] ^ m[268] ^ m[270] ^ m[273] ^ m[275] ^ m[277] ^ m[279] ^ m[281] ^ m[283] ^ m[285] ^ m[287] ^ m[289] ^ m[291] ^ m[293] ^ m[295] ^ m[297] ^ m[299] ^ m[301] ^ m[303] ^ m[305] ^ m[307] ^ m[309] ^ m[311] ^ m[313] ^ m[315] ^ m[317] ^ m[319] ^ m[321] ^ m[323] ^ m[325] ^ m[327] ^ m[329] ^ m[331] ^ m[333] ^ m[335] ^ m[337] ^ m[339] ^ m[341] ^ m[343] ^ m[345] ^ m[347] ^ m[349] ^ m[351] ^ m[353] ^ m[355] ^ m[357] ^ m[359] ^ m[361] ^ m[363] ^ m[365] ^ m[367] ^ m[369] ^ m[371] ^ m[373] ^ m[375] ^ m[377] ^ m[379] ^ m[381] ^ m[383] ^ m[385] ^ m[387] ^ m[389] ^ m[391] ^ m[393] ^ m[395] ^ m[397] ^ m[399] ^ m[401] ^ m[403] ^ m[405] ^ m[407] ^ m[409] ^ m[411] ^ m[413] ^ m[415] ^ m[417] ^ m[419] ^ m[421] ^ m[423] ^ m[425] ^ m[427] ^ m[429] ^ m[431] ^ m[433] ^ m[435] ^ m[437] ^ m[439] ^ m[440] ^ m[442] ^ m[444] ^ m[446] ^ m[448] ^ m[450] ^ m[452] ^ m[454] ^ m[456] ^ m[458] ^ m[460] ^ m[462] ^ m[464] ^ m[466] ^ m[468] ^ m[470] ^ m[472] ^ m[474] ^ m[476] ^ m[478] ^ m[480] ^ m[482] ^ m[484] ^ m[486] ^ m[488] ^ m[490] ^ m[492] ^ m[494] ^ m[496] ^ m[498] ^ m[500] ^ m[502] ^ m[504] ^ m[506] ^ m[508] ^ m[510] ^ m[513] ^ m[515] ^ m[517] ^ m[519] ^ m[521] ^ m[523] ^ m[525] ^ m[527] ^ m[529] ^ m[531] ^ m[533] ^ m[535] ^ m[537] ^ m[539] ^ m[541] ^ m[543] ^ m[545] ^ m[547] ^ m[549] ^ m[551] ^ m[553] ^ m[555] ^ m[557] ^ m[559] ^ m[561] ^ m[563] ^ m[565] ^ m[567] ^ m[569] ^ m[571] ^ m[573] ^ m[575] ^ m[577] ^ m[579] ^ m[581] ^ m[583] ^ m[585] ^ m[587] ^ m[589] ^ m[591] ^ m[593] ^ m[595] ^ m[597] ^ m[599] ^ m[601] ^ m[603] ^ m[605] ^ m[607] ^ m[609] ^ m[611] ^ m[613] ^ m[615] ^ m[617] ^ m[619] ^ m[621] ^ m[623] ^ m[625] ^ m[627] ^ m[629] ^ m[631] ^ m[633] ^ m[635] ^ m[637] ^ m[639] ^ m[641] ^ m[643] ^ m[645] ^ m[647] ^ m[649] ^ m[651] ^ m[653] ^ m[655] ^ m[657] ^ m[659] ^ m[661] ^ m[663] ^ m[665] ^ m[667] ^ m[669] ^ m[671] ^ m[673] ^ m[675] ^ m[677] ^ m[679] ^ m[680] ^ m[682] ^ m[684] ^ m[686] ^ m[688] ^ m[690] ^ m[692] ^ m[694] ^ m[696] ^ m[698] ^ m[700] ^ m[702] ^ m[704] ^ m[706] ^ m[708] ^ m[710] ^ m[712] ^ m[714] ^ m[716] ^ m[718] ^ m[720] ^ m[722] ^ m[724] ^ m[726] ^ m[728] ^ m[730] ^ m[732] ^ m[734] ^ m[736] ^ m[738] ^ m[740] ^ m[742] ^ m[744] ^ m[746] ^ m[748] ^ m[750] ^ m[752] ^ m[754] ^ m[756] ^ m[758] ^ m[760] ^ m[762] ^ m[764] ^ m[766] ^ m[768] ^ m[770] ^ m[772] ^ m[774] ^ m[776] ^ m[778] ^ m[780] ^ m[782] ^ m[784] ^ m[786] ^ m[788] ^ m[790] ^ m[792] ^ m[794] ^ m[796] ^ m[798] ^ m[800] ^ m[802] ^ m[804] ^ m[806] ^ m[808] ^ m[810] ^ m[812] ^ m[814] ^ m[816] ^ m[818] ^ m[820] ^ m[822] ^ m[824] ^ m[826] ^ m[828] ^ m[830] ^ m[832] ^ m[834] ^ m[836] ^ m[838] ^ m[840] ^ m[842] ^ m[844] ^ m[846] ^ m[849] ^ m[851] ^ m[853] ^ m[855] ^ m[857] ^ m[859] ^ m[861] ^ m[863] ^ m[865] ^ m[867] ^ m[869] ^ m[871] ^ m[873] ^ m[875] ^ m[877] ^ m[879] ^ m[881] ^ m[883] ^ m[885] ^ m[887] ^ m[889] ^ m[891] ^ m[893] ^ m[895] ^ m[897] ^ m[899] ^ m[901] ^ m[903] ^ m[905] ^ m[907] ^ m[909] ^ m[911] ^ m[913] ^ m[915] ^ m[917] ^ m[919] ^ m[921] ^ m[923] ^ m[925] ^ m[927] ^ m[929] ^ m[931] ^ m[933] ^ m[935] ^ m[937] ^ m[939] ^ m[941] ^ m[943] ^ m[945] ^ m[947] ^ m[949] ^ m[951] ^ m[953] ^ m[955] ^ m[957] ^ m[959] ^ m[961] ^ m[963] ^ m[965] ^ m[967] ^ m[969] ^ m[971] ^ m[973] ^ m[975] ^ m[977] ^ m[979] ^ m[981] ^ m[983] ^ m[985] ^ m[987] ^ m[989] ^ m[991] ^ m[993] ^ m[995] ^ m[997] ^ m[999] ^ m[1001] ^ m[1003] ^ m[1005] ^ m[1007] ^ m[1009] ^ m[1011] ^ m[1013] ^ m[1015] ^ m[1017] ^ m[1019] ^ m[1021] ^ m[1023] ^ m[1025] ^ m[1027] ^ m[1029] ^ m[1031] ^ m[1033] ^ m[1035] ^ m[1037] ^ m[1039] ^ m[1041] ^ m[1043] ^ m[1045] ^ m[1047] ^ m[1049] ^ m[1051] ^ m[1053] ^ m[1055] ^ m[1057] ^ m[1059] ^ m[1061] ^ m[1063] ^ m[1065] ^ m[1067] ^ m[1069] ^ m[1071] ^ m[1073] ^ m[1075] ^ m[1077] ^ m[1079] ^ m[1081] ^ m[1083] ^ m[1085] ^ m[1087] ^ m[1089] ^ m[1091] ^ m[1093] ^ m[1095] ^ m[1097] ^ m[1099] ^ m[1100] ^ m[1102] ^ m[1104] ^ m[1106] ^ m[1108] ^ m[1110] ^ m[1112] ^ m[1114] ^ m[1116] ^ m[1118] ^ m[1120] ^ m[1122] ^ m[1124] ^ m[1126] ^ m[1128] ^ m[1130] ^ m[1132] ^ m[1134] ^ m[1136] ^ m[1138] ^ m[1140] ^ m[1142] ^ m[1144] ^ m[1146] ^ m[1148] ^ m[1150] ^ m[1152] ^ m[1154] ^ m[1156] ^ m[1158] ^ m[1160] ^ m[1162] ^ m[1164] ^ m[1166] ^ m[1168] ^ m[1170] ^ m[1172] ^ m[1174] ^ m[1176] ^ m[1178] ^ m[1180] ^ m[1182] ^ m[1184] ^ m[1186] ^ m[1188] ^ m[1190] ^ m[1192] ^ m[1194] ^ m[1196] ^ m[1198] ^ m[1200] ^ m[1202] ^ m[1204] ^ m[1206] ^ m[1208] ^ m[1210] ^ m[1212] ^ m[1214] ^ m[1216] ^ m[1218] ^ m[1220] ^ m[1222] ^ m[1224] ^ m[1226] ^ m[1228] ^ m[1230] ^ m[1232] ^ m[1234] ^ m[1236] ^ m[1238] ^ m[1240] ^ m[1242] ^ m[1244] ^ m[1246] ^ m[1248] ^ m[1250] ^ m[1252] ^ m[1254] ^ m[1256] ^ m[1258] ^ m[1260] ^ m[1262] ^ m[1264] ^ m[1266] ^ m[1269] ^ m[1271] ^ m[1273] ^ m[1275] ^ m[1277] ^ m[1279] ^ m[1281] ^ m[1283] ^ m[1285] ^ m[1287] ^ m[1289] ^ m[1291] ^ m[1293] ^ m[1295] ^ m[1297] ^ m[1299] ^ m[1301] ^ m[1303] ^ m[1305] ^ m[1307] ^ m[1309] ^ m[1311] ^ m[1313] ^ m[1315] ^ m[1317] ^ m[1319] ^ m[1321] ^ m[1323] ^ m[1325] ^ m[1327] ^ m[1329] ^ m[1331] ^ m[1333] ^ m[1335] ^ m[1337] ^ m[1339] ^ m[1341] ^ m[1343] ^ m[1345] ^ m[1347] ^ m[1349] ^ m[1351] ^ m[1353] ^ m[1355] ^ m[1357] ^ m[1359] ^ m[1361] ^ m[1363] ^ m[1365] ^ m[1367] ^ m[1369] ^ m[1371] ^ m[1373] ^ m[1375] ^ m[1377] ^ m[1379] ^ m[1381] ^ m[1383] ^ m[1385] ^ m[1387] ^ m[1389] ^ m[1391] ^ m[1393] ^ m[1395] ^ m[1397] ^ m[1399] ^ m[1401] ^ m[1403] ^ m[1405] ^ m[1407] ^ m[1409] ^ m[1411] ^ m[1413] ^ m[1415] ^ m[1417] ^ m[1419] ^ m[1421] ^ m[1423] ^ m[1425] ^ m[1427] ^ m[1429] ^ m[1431] ^ m[1433] ^ m[1435] ^ m[1437] ^ m[1439] ^ m[1441] ^ m[1443] ^ m[1445] ^ m[1447] ^ m[1449] ^ m[1451] ^ m[1453] ^ m[1455] ^ m[1457] ^ m[1459] ^ m[1461] ^ m[1463] ^ m[1465] ^ m[1467] ^ m[1469] ^ m[1471] ^ m[1473] ^ m[1475] ^ m[1477] ^ m[1479] ^ m[1481] ^ m[1483] ^ m[1485] ^ m[1487] ^ m[1489] ^ m[1491] ^ m[1493] ^ m[1495] ^ m[1497] ^ m[1499] ^ m[1501] ^ m[1503] ^ m[1505] ^ m[1507] ^ m[1509] ^ m[1511] ^ m[1513] ^ m[1515] ^ m[1517] ^ m[1519] ^ m[1520] ^ m[1522] ^ m[1524] ^ m[1526] ^ m[1528] ^ m[1530] ^ m[1532] ^ m[1534] ^ m[1536] ^ m[1538] ^ m[1540] ^ m[1542] ^ m[1544] ^ m[1546] ^ m[1548] ^ m[1550] ^ m[1552] ^ m[1554] ^ m[1556] ^ m[1558] ^ m[1560] ^ m[1562] ^ m[1564] ^ m[1566] ^ m[1568] ^ m[1570] ^ m[1572] ^ m[1574] ^ m[1576] ^ m[1578] ^ m[1580] ^ m[1582] ^ m[1584] ^ m[1586] ^ m[1588] ^ m[1590] ^ m[1592] ^ m[1594] ^ m[1596] ^ m[1598] ^ m[1600] ^ m[1602] ^ m[1604] ^ m[1606] ^ m[1608] ^ m[1610] ^ m[1612] ^ m[1614] ^ m[1616] ^ m[1618] ^ m[1620] ^ m[1622] ^ m[1624] ^ m[1626] ^ m[1628] ^ m[1630] ^ m[1632] ^ m[1634] ^ m[1636] ^ m[1638] ^ m[1640] ^ m[1642] ^ m[1644] ^ m[1646] ^ m[1648] ^ m[1650] ^ m[1652] ^ m[1654] ^ m[1656] ^ m[1658] ^ m[1660] ^ m[1662] ^ m[1664] ^ m[1666] ^ m[1668] ^ m[1670] ^ m[1672] ^ m[1674] ^ m[1676] ^ m[1678] ^ m[1680] ^ m[1682] ^ m[1684] ^ m[1686] ^ m[1688] ^ m[1690] ^ m[1692] ^ m[1694] ^ m[1696] ^ m[1698] ^ m[1700] ^ m[1702] ^ m[1704] ^ m[1706] ^ m[1708] ^ m[1710] ^ m[1712] ^ m[1714] ^ m[1716] ^ m[1718] ^ m[1720] ^ m[1722] ^ m[1724] ^ m[1726] ^ m[1728] ^ m[1730] ^ m[1732] ^ m[1734] ^ m[1736] ^ m[1738] ^ m[1740] ^ m[1742] ^ m[1744] ^ m[1746] ^ m[1748] ^ m[1750] ^ m[1752] ^ m[1754] ^ m[1756] ^ m[1758] ^ m[1760] ^ m[1762] ^ m[1764] ^ m[1766] ^ m[1768] ^ m[1770] ^ m[1773] ^ m[1775] ^ m[1777] ^ m[1779] ^ m[1781] ^ m[1783] ^ m[1785] ^ m[1787] ^ m[1789] ^ m[1791] ^ m[1793] ^ m[1795] ^ m[1797] ^ m[1799] ^ m[1801] ^ m[1803] ^ m[1805] ^ m[1807] ^ m[1809] ^ m[1811] ^ m[1813] ^ m[1815] ^ m[1817] ^ m[1819] ^ m[1821] ^ m[1823] ^ m[1825] ^ m[1827] ^ m[1829] ^ m[1831] ^ m[1833] ^ m[1835] ^ m[1837] ^ m[1839] ^ m[1841] ^ m[1843] ^ m[1845] ^ m[1847] ^ m[1849] ^ m[1851] ^ m[1853] ^ m[1855] ^ m[1857] ^ m[1859] ^ m[1861] ^ m[1863] ^ m[1865] ^ m[1867] ^ m[1869] ^ m[1871] ^ m[1873] ^ m[1875] ^ m[1877] ^ m[1879] ^ m[1881] ^ m[1883] ^ m[1885] ^ m[1887] ^ m[1889] ^ m[1891] ^ m[1893] ^ m[1895] ^ m[1897] ^ m[1899] ^ m[1901] ^ m[1903] ^ m[1905] ^ m[1907] ^ m[1909] ^ m[1911] ^ m[1913] ^ m[1915] ^ m[1917] ^ m[1919] ^ m[1921] ^ m[1923] ^ m[1925] ^ m[1927] ^ m[1929] ^ m[1931] ^ m[1933] ^ m[1935] ^ m[1937] ^ m[1939] ^ m[1941] ^ m[1943] ^ m[1945] ^ m[1947] ^ m[1949] ^ m[1951] ^ m[1953] ^ m[1955] ^ m[1957] ^ m[1959] ^ m[1961] ^ m[1963] ^ m[1965] ^ m[1967] ^ m[1969] ^ m[1971] ^ m[1973] ^ m[1975] ^ m[1977] ^ m[1979] ^ m[1981] ^ m[1983] ^ m[1985] ^ m[1987] ^ m[1989] ^ m[1991] ^ m[1993] ^ m[1995] ^ m[1997] ^ m[1999] ^ m[2001] ^ m[2003] ^ m[2005] ^ m[2007] ^ m[2009] ^ m[2011] ^ m[2013] ^ m[2015] ^ m[2017] ^ m[2019] ^ m[2021] ^ m[2023] ^ m[2024] ^ m[2025] ^ m[2026] ^ m[2027] ^ m[2028] ^ m[2029] ^ m[2030] ^ m[2031] ^ m[2032] ^ m[2034] ^ m[2035];
    assign parity[10] = m[0] ^ m[2] ^ m[4] ^ m[6] ^ m[8] ^ m[10] ^ m[12] ^ m[14] ^ m[16] ^ m[18] ^ m[21] ^ m[23] ^ m[25] ^ m[27] ^ m[29] ^ m[31] ^ m[33] ^ m[35] ^ m[37] ^ m[39] ^ m[41] ^ m[43] ^ m[45] ^ m[47] ^ m[49] ^ m[51] ^ m[53] ^ m[55] ^ m[57] ^ m[59] ^ m[61] ^ m[63] ^ m[65] ^ m[67] ^ m[69] ^ m[71] ^ m[73] ^ m[75] ^ m[77] ^ m[79] ^ m[81] ^ m[83] ^ m[85] ^ m[87] ^ m[89] ^ m[91] ^ m[93] ^ m[95] ^ m[97] ^ m[99] ^ m[101] ^ m[103] ^ m[105] ^ m[107] ^ m[109] ^ m[110] ^ m[112] ^ m[114] ^ m[116] ^ m[118] ^ m[120] ^ m[122] ^ m[124] ^ m[126] ^ m[128] ^ m[130] ^ m[132] ^ m[134] ^ m[136] ^ m[138] ^ m[140] ^ m[142] ^ m[144] ^ m[146] ^ m[148] ^ m[150] ^ m[152] ^ m[154] ^ m[156] ^ m[158] ^ m[160] ^ m[162] ^ m[164] ^ m[166] ^ m[168] ^ m[170] ^ m[172] ^ m[174] ^ m[176] ^ m[178] ^ m[180] ^ m[182] ^ m[184] ^ m[186] ^ m[188] ^ m[190] ^ m[192] ^ m[194] ^ m[196] ^ m[198] ^ m[201] ^ m[203] ^ m[205] ^ m[207] ^ m[209] ^ m[211] ^ m[213] ^ m[215] ^ m[217] ^ m[219] ^ m[221] ^ m[223] ^ m[225] ^ m[227] ^ m[229] ^ m[231] ^ m[233] ^ m[235] ^ m[237] ^ m[239] ^ m[241] ^ m[243] ^ m[245] ^ m[247] ^ m[249] ^ m[251] ^ m[253] ^ m[255] ^ m[257] ^ m[259] ^ m[261] ^ m[263] ^ m[265] ^ m[267] ^ m[269] ^ m[271] ^ m[273] ^ m[275] ^ m[277] ^ m[279] ^ m[281] ^ m[283] ^ m[285] ^ m[287] ^ m[289] ^ m[291] ^ m[293] ^ m[295] ^ m[297] ^ m[299] ^ m[301] ^ m[303] ^ m[305] ^ m[307] ^ m[309] ^ m[311] ^ m[313] ^ m[315] ^ m[317] ^ m[319] ^ m[321] ^ m[323] ^ m[325] ^ m[327] ^ m[329] ^ m[331] ^ m[333] ^ m[335] ^ m[337] ^ m[339] ^ m[341] ^ m[343] ^ m[345] ^ m[347] ^ m[349] ^ m[351] ^ m[353] ^ m[355] ^ m[357] ^ m[359] ^ m[361] ^ m[363] ^ m[365] ^ m[367] ^ m[369] ^ m[371] ^ m[373] ^ m[375] ^ m[377] ^ m[379] ^ m[381] ^ m[383] ^ m[385] ^ m[387] ^ m[389] ^ m[391] ^ m[393] ^ m[395] ^ m[397] ^ m[399] ^ m[401] ^ m[403] ^ m[405] ^ m[407] ^ m[409] ^ m[411] ^ m[413] ^ m[415] ^ m[417] ^ m[419] ^ m[421] ^ m[423] ^ m[425] ^ m[427] ^ m[429] ^ m[431] ^ m[433] ^ m[435] ^ m[437] ^ m[439] ^ m[440] ^ m[442] ^ m[444] ^ m[446] ^ m[448] ^ m[450] ^ m[452] ^ m[454] ^ m[456] ^ m[458] ^ m[460] ^ m[462] ^ m[464] ^ m[466] ^ m[468] ^ m[470] ^ m[472] ^ m[474] ^ m[476] ^ m[478] ^ m[480] ^ m[482] ^ m[484] ^ m[486] ^ m[488] ^ m[490] ^ m[492] ^ m[494] ^ m[496] ^ m[498] ^ m[500] ^ m[502] ^ m[504] ^ m[506] ^ m[508] ^ m[510] ^ m[512] ^ m[514] ^ m[516] ^ m[518] ^ m[520] ^ m[522] ^ m[524] ^ m[526] ^ m[528] ^ m[530] ^ m[532] ^ m[534] ^ m[536] ^ m[538] ^ m[540] ^ m[542] ^ m[544] ^ m[546] ^ m[548] ^ m[550] ^ m[552] ^ m[554] ^ m[556] ^ m[558] ^ m[560] ^ m[562] ^ m[564] ^ m[566] ^ m[568] ^ m[570] ^ m[572] ^ m[574] ^ m[576] ^ m[578] ^ m[580] ^ m[582] ^ m[584] ^ m[586] ^ m[588] ^ m[590] ^ m[592] ^ m[594] ^ m[596] ^ m[598] ^ m[600] ^ m[602] ^ m[604] ^ m[606] ^ m[608] ^ m[610] ^ m[612] ^ m[614] ^ m[616] ^ m[618] ^ m[620] ^ m[622] ^ m[624] ^ m[626] ^ m[628] ^ m[630] ^ m[632] ^ m[634] ^ m[636] ^ m[638] ^ m[640] ^ m[642] ^ m[644] ^ m[646] ^ m[648] ^ m[650] ^ m[652] ^ m[654] ^ m[656] ^ m[658] ^ m[660] ^ m[662] ^ m[664] ^ m[666] ^ m[668] ^ m[670] ^ m[672] ^ m[674] ^ m[676] ^ m[678] ^ m[681] ^ m[683] ^ m[685] ^ m[687] ^ m[689] ^ m[691] ^ m[693] ^ m[695] ^ m[697] ^ m[699] ^ m[701] ^ m[703] ^ m[705] ^ m[707] ^ m[709] ^ m[711] ^ m[713] ^ m[715] ^ m[717] ^ m[719] ^ m[721] ^ m[723] ^ m[725] ^ m[727] ^ m[729] ^ m[731] ^ m[733] ^ m[735] ^ m[737] ^ m[739] ^ m[741] ^ m[743] ^ m[745] ^ m[747] ^ m[749] ^ m[751] ^ m[753] ^ m[755] ^ m[757] ^ m[759] ^ m[761] ^ m[763] ^ m[765] ^ m[767] ^ m[769] ^ m[771] ^ m[773] ^ m[775] ^ m[777] ^ m[779] ^ m[781] ^ m[783] ^ m[785] ^ m[787] ^ m[789] ^ m[791] ^ m[793] ^ m[795] ^ m[797] ^ m[799] ^ m[801] ^ m[803] ^ m[805] ^ m[807] ^ m[809] ^ m[811] ^ m[813] ^ m[815] ^ m[817] ^ m[819] ^ m[821] ^ m[823] ^ m[825] ^ m[827] ^ m[829] ^ m[831] ^ m[833] ^ m[835] ^ m[837] ^ m[839] ^ m[841] ^ m[843] ^ m[845] ^ m[847] ^ m[849] ^ m[851] ^ m[853] ^ m[855] ^ m[857] ^ m[859] ^ m[861] ^ m[863] ^ m[865] ^ m[867] ^ m[869] ^ m[871] ^ m[873] ^ m[875] ^ m[877] ^ m[879] ^ m[881] ^ m[883] ^ m[885] ^ m[887] ^ m[889] ^ m[891] ^ m[893] ^ m[895] ^ m[897] ^ m[899] ^ m[901] ^ m[903] ^ m[905] ^ m[907] ^ m[909] ^ m[911] ^ m[913] ^ m[915] ^ m[917] ^ m[919] ^ m[921] ^ m[923] ^ m[925] ^ m[927] ^ m[929] ^ m[931] ^ m[933] ^ m[935] ^ m[937] ^ m[939] ^ m[941] ^ m[943] ^ m[945] ^ m[947] ^ m[949] ^ m[951] ^ m[953] ^ m[955] ^ m[957] ^ m[959] ^ m[961] ^ m[963] ^ m[965] ^ m[967] ^ m[969] ^ m[971] ^ m[973] ^ m[975] ^ m[977] ^ m[979] ^ m[981] ^ m[983] ^ m[985] ^ m[987] ^ m[989] ^ m[991] ^ m[993] ^ m[995] ^ m[997] ^ m[999] ^ m[1001] ^ m[1003] ^ m[1005] ^ m[1007] ^ m[1009] ^ m[1011] ^ m[1013] ^ m[1015] ^ m[1017] ^ m[1019] ^ m[1021] ^ m[1023] ^ m[1025] ^ m[1027] ^ m[1029] ^ m[1031] ^ m[1033] ^ m[1035] ^ m[1037] ^ m[1039] ^ m[1041] ^ m[1043] ^ m[1045] ^ m[1047] ^ m[1049] ^ m[1051] ^ m[1053] ^ m[1055] ^ m[1057] ^ m[1059] ^ m[1061] ^ m[1063] ^ m[1065] ^ m[1067] ^ m[1069] ^ m[1071] ^ m[1073] ^ m[1075] ^ m[1077] ^ m[1079] ^ m[1081] ^ m[1083] ^ m[1085] ^ m[1087] ^ m[1089] ^ m[1091] ^ m[1093] ^ m[1095] ^ m[1097] ^ m[1099] ^ m[1100] ^ m[1102] ^ m[1104] ^ m[1106] ^ m[1108] ^ m[1110] ^ m[1112] ^ m[1114] ^ m[1116] ^ m[1118] ^ m[1120] ^ m[1122] ^ m[1124] ^ m[1126] ^ m[1128] ^ m[1130] ^ m[1132] ^ m[1134] ^ m[1136] ^ m[1138] ^ m[1140] ^ m[1142] ^ m[1144] ^ m[1146] ^ m[1148] ^ m[1150] ^ m[1152] ^ m[1154] ^ m[1156] ^ m[1158] ^ m[1160] ^ m[1162] ^ m[1164] ^ m[1166] ^ m[1168] ^ m[1170] ^ m[1172] ^ m[1174] ^ m[1176] ^ m[1178] ^ m[1180] ^ m[1182] ^ m[1184] ^ m[1186] ^ m[1188] ^ m[1190] ^ m[1192] ^ m[1194] ^ m[1196] ^ m[1198] ^ m[1200] ^ m[1202] ^ m[1204] ^ m[1206] ^ m[1208] ^ m[1210] ^ m[1212] ^ m[1214] ^ m[1216] ^ m[1218] ^ m[1220] ^ m[1222] ^ m[1224] ^ m[1226] ^ m[1228] ^ m[1230] ^ m[1232] ^ m[1234] ^ m[1236] ^ m[1238] ^ m[1240] ^ m[1242] ^ m[1244] ^ m[1246] ^ m[1248] ^ m[1250] ^ m[1252] ^ m[1254] ^ m[1256] ^ m[1258] ^ m[1260] ^ m[1262] ^ m[1264] ^ m[1266] ^ m[1268] ^ m[1270] ^ m[1272] ^ m[1274] ^ m[1276] ^ m[1278] ^ m[1280] ^ m[1282] ^ m[1284] ^ m[1286] ^ m[1288] ^ m[1290] ^ m[1292] ^ m[1294] ^ m[1296] ^ m[1298] ^ m[1300] ^ m[1302] ^ m[1304] ^ m[1306] ^ m[1308] ^ m[1310] ^ m[1312] ^ m[1314] ^ m[1316] ^ m[1318] ^ m[1320] ^ m[1322] ^ m[1324] ^ m[1326] ^ m[1328] ^ m[1330] ^ m[1332] ^ m[1334] ^ m[1336] ^ m[1338] ^ m[1340] ^ m[1342] ^ m[1344] ^ m[1346] ^ m[1348] ^ m[1350] ^ m[1352] ^ m[1354] ^ m[1356] ^ m[1358] ^ m[1360] ^ m[1362] ^ m[1364] ^ m[1366] ^ m[1368] ^ m[1370] ^ m[1372] ^ m[1374] ^ m[1376] ^ m[1378] ^ m[1380] ^ m[1382] ^ m[1384] ^ m[1386] ^ m[1388] ^ m[1390] ^ m[1392] ^ m[1394] ^ m[1396] ^ m[1398] ^ m[1400] ^ m[1402] ^ m[1404] ^ m[1406] ^ m[1408] ^ m[1410] ^ m[1412] ^ m[1414] ^ m[1416] ^ m[1418] ^ m[1420] ^ m[1422] ^ m[1424] ^ m[1426] ^ m[1428] ^ m[1430] ^ m[1432] ^ m[1434] ^ m[1436] ^ m[1438] ^ m[1440] ^ m[1442] ^ m[1444] ^ m[1446] ^ m[1448] ^ m[1450] ^ m[1452] ^ m[1454] ^ m[1456] ^ m[1458] ^ m[1460] ^ m[1462] ^ m[1464] ^ m[1466] ^ m[1468] ^ m[1470] ^ m[1472] ^ m[1474] ^ m[1476] ^ m[1478] ^ m[1480] ^ m[1482] ^ m[1484] ^ m[1486] ^ m[1488] ^ m[1490] ^ m[1492] ^ m[1494] ^ m[1496] ^ m[1498] ^ m[1500] ^ m[1502] ^ m[1504] ^ m[1506] ^ m[1508] ^ m[1510] ^ m[1512] ^ m[1514] ^ m[1516] ^ m[1518] ^ m[1521] ^ m[1523] ^ m[1525] ^ m[1527] ^ m[1529] ^ m[1531] ^ m[1533] ^ m[1535] ^ m[1537] ^ m[1539] ^ m[1541] ^ m[1543] ^ m[1545] ^ m[1547] ^ m[1549] ^ m[1551] ^ m[1553] ^ m[1555] ^ m[1557] ^ m[1559] ^ m[1561] ^ m[1563] ^ m[1565] ^ m[1567] ^ m[1569] ^ m[1571] ^ m[1573] ^ m[1575] ^ m[1577] ^ m[1579] ^ m[1581] ^ m[1583] ^ m[1585] ^ m[1587] ^ m[1589] ^ m[1591] ^ m[1593] ^ m[1595] ^ m[1597] ^ m[1599] ^ m[1601] ^ m[1603] ^ m[1605] ^ m[1607] ^ m[1609] ^ m[1611] ^ m[1613] ^ m[1615] ^ m[1617] ^ m[1619] ^ m[1621] ^ m[1623] ^ m[1625] ^ m[1627] ^ m[1629] ^ m[1631] ^ m[1633] ^ m[1635] ^ m[1637] ^ m[1639] ^ m[1641] ^ m[1643] ^ m[1645] ^ m[1647] ^ m[1649] ^ m[1651] ^ m[1653] ^ m[1655] ^ m[1657] ^ m[1659] ^ m[1661] ^ m[1663] ^ m[1665] ^ m[1667] ^ m[1669] ^ m[1671] ^ m[1673] ^ m[1675] ^ m[1677] ^ m[1679] ^ m[1681] ^ m[1683] ^ m[1685] ^ m[1687] ^ m[1689] ^ m[1691] ^ m[1693] ^ m[1695] ^ m[1697] ^ m[1699] ^ m[1701] ^ m[1703] ^ m[1705] ^ m[1707] ^ m[1709] ^ m[1711] ^ m[1713] ^ m[1715] ^ m[1717] ^ m[1719] ^ m[1721] ^ m[1723] ^ m[1725] ^ m[1727] ^ m[1729] ^ m[1731] ^ m[1733] ^ m[1735] ^ m[1737] ^ m[1739] ^ m[1741] ^ m[1743] ^ m[1745] ^ m[1747] ^ m[1749] ^ m[1751] ^ m[1753] ^ m[1755] ^ m[1757] ^ m[1759] ^ m[1761] ^ m[1763] ^ m[1765] ^ m[1767] ^ m[1769] ^ m[1771] ^ m[1773] ^ m[1775] ^ m[1777] ^ m[1779] ^ m[1781] ^ m[1783] ^ m[1785] ^ m[1787] ^ m[1789] ^ m[1791] ^ m[1793] ^ m[1795] ^ m[1797] ^ m[1799] ^ m[1801] ^ m[1803] ^ m[1805] ^ m[1807] ^ m[1809] ^ m[1811] ^ m[1813] ^ m[1815] ^ m[1817] ^ m[1819] ^ m[1821] ^ m[1823] ^ m[1825] ^ m[1827] ^ m[1829] ^ m[1831] ^ m[1833] ^ m[1835] ^ m[1837] ^ m[1839] ^ m[1841] ^ m[1843] ^ m[1845] ^ m[1847] ^ m[1849] ^ m[1851] ^ m[1853] ^ m[1855] ^ m[1857] ^ m[1859] ^ m[1861] ^ m[1863] ^ m[1865] ^ m[1867] ^ m[1869] ^ m[1871] ^ m[1873] ^ m[1875] ^ m[1877] ^ m[1879] ^ m[1881] ^ m[1883] ^ m[1885] ^ m[1887] ^ m[1889] ^ m[1891] ^ m[1893] ^ m[1895] ^ m[1897] ^ m[1899] ^ m[1901] ^ m[1903] ^ m[1905] ^ m[1907] ^ m[1909] ^ m[1911] ^ m[1913] ^ m[1915] ^ m[1917] ^ m[1919] ^ m[1921] ^ m[1923] ^ m[1925] ^ m[1927] ^ m[1929] ^ m[1931] ^ m[1933] ^ m[1935] ^ m[1937] ^ m[1939] ^ m[1941] ^ m[1943] ^ m[1945] ^ m[1947] ^ m[1949] ^ m[1951] ^ m[1953] ^ m[1955] ^ m[1957] ^ m[1959] ^ m[1961] ^ m[1963] ^ m[1965] ^ m[1967] ^ m[1969] ^ m[1971] ^ m[1973] ^ m[1975] ^ m[1977] ^ m[1979] ^ m[1981] ^ m[1983] ^ m[1985] ^ m[1987] ^ m[1989] ^ m[1991] ^ m[1993] ^ m[1995] ^ m[1997] ^ m[1999] ^ m[2001] ^ m[2003] ^ m[2005] ^ m[2007] ^ m[2009] ^ m[2011] ^ m[2013] ^ m[2015] ^ m[2017] ^ m[2019] ^ m[2021] ^ m[2023] ^ m[2024] ^ m[2025] ^ m[2026] ^ m[2027] ^ m[2028] ^ m[2029] ^ m[2030] ^ m[2031] ^ m[2032] ^ m[2033] ^ m[2035];
    assign parity[11] = m[0] ^ m[2] ^ m[4] ^ m[6] ^ m[8] ^ m[10] ^ m[12] ^ m[14] ^ m[16] ^ m[18] ^ m[20] ^ m[22] ^ m[24] ^ m[26] ^ m[28] ^ m[30] ^ m[32] ^ m[34] ^ m[36] ^ m[38] ^ m[40] ^ m[42] ^ m[44] ^ m[46] ^ m[48] ^ m[50] ^ m[52] ^ m[54] ^ m[56] ^ m[58] ^ m[60] ^ m[62] ^ m[64] ^ m[66] ^ m[68] ^ m[70] ^ m[72] ^ m[74] ^ m[76] ^ m[78] ^ m[80] ^ m[82] ^ m[84] ^ m[86] ^ m[88] ^ m[90] ^ m[92] ^ m[94] ^ m[96] ^ m[98] ^ m[100] ^ m[102] ^ m[104] ^ m[106] ^ m[108] ^ m[111] ^ m[113] ^ m[115] ^ m[117] ^ m[119] ^ m[121] ^ m[123] ^ m[125] ^ m[127] ^ m[129] ^ m[131] ^ m[133] ^ m[135] ^ m[137] ^ m[139] ^ m[141] ^ m[143] ^ m[145] ^ m[147] ^ m[149] ^ m[151] ^ m[153] ^ m[155] ^ m[157] ^ m[159] ^ m[161] ^ m[163] ^ m[165] ^ m[167] ^ m[169] ^ m[171] ^ m[173] ^ m[175] ^ m[177] ^ m[179] ^ m[181] ^ m[183] ^ m[185] ^ m[187] ^ m[189] ^ m[191] ^ m[193] ^ m[195] ^ m[197] ^ m[199] ^ m[201] ^ m[203] ^ m[205] ^ m[207] ^ m[209] ^ m[211] ^ m[213] ^ m[215] ^ m[217] ^ m[219] ^ m[221] ^ m[223] ^ m[225] ^ m[227] ^ m[229] ^ m[231] ^ m[233] ^ m[235] ^ m[237] ^ m[239] ^ m[241] ^ m[243] ^ m[245] ^ m[247] ^ m[249] ^ m[251] ^ m[253] ^ m[255] ^ m[257] ^ m[259] ^ m[261] ^ m[263] ^ m[265] ^ m[267] ^ m[269] ^ m[271] ^ m[273] ^ m[275] ^ m[277] ^ m[279] ^ m[281] ^ m[283] ^ m[285] ^ m[287] ^ m[289] ^ m[291] ^ m[293] ^ m[295] ^ m[297] ^ m[299] ^ m[301] ^ m[303] ^ m[305] ^ m[307] ^ m[309] ^ m[311] ^ m[313] ^ m[315] ^ m[317] ^ m[319] ^ m[321] ^ m[323] ^ m[325] ^ m[327] ^ m[329] ^ m[331] ^ m[333] ^ m[335] ^ m[337] ^ m[339] ^ m[341] ^ m[343] ^ m[345] ^ m[347] ^ m[349] ^ m[351] ^ m[353] ^ m[355] ^ m[357] ^ m[359] ^ m[361] ^ m[363] ^ m[365] ^ m[367] ^ m[369] ^ m[371] ^ m[373] ^ m[375] ^ m[377] ^ m[379] ^ m[381] ^ m[383] ^ m[385] ^ m[387] ^ m[389] ^ m[391] ^ m[393] ^ m[395] ^ m[397] ^ m[399] ^ m[401] ^ m[403] ^ m[405] ^ m[407] ^ m[409] ^ m[411] ^ m[413] ^ m[415] ^ m[417] ^ m[419] ^ m[421] ^ m[423] ^ m[425] ^ m[427] ^ m[429] ^ m[431] ^ m[433] ^ m[435] ^ m[437] ^ m[439] ^ m[440] ^ m[442] ^ m[444] ^ m[446] ^ m[448] ^ m[450] ^ m[452] ^ m[454] ^ m[456] ^ m[458] ^ m[460] ^ m[462] ^ m[464] ^ m[466] ^ m[468] ^ m[470] ^ m[472] ^ m[474] ^ m[476] ^ m[478] ^ m[480] ^ m[482] ^ m[484] ^ m[486] ^ m[488] ^ m[490] ^ m[492] ^ m[494] ^ m[496] ^ m[498] ^ m[500] ^ m[502] ^ m[504] ^ m[506] ^ m[508] ^ m[510] ^ m[512] ^ m[514] ^ m[516] ^ m[518] ^ m[520] ^ m[522] ^ m[524] ^ m[526] ^ m[528] ^ m[530] ^ m[532] ^ m[534] ^ m[536] ^ m[538] ^ m[540] ^ m[542] ^ m[544] ^ m[546] ^ m[548] ^ m[550] ^ m[552] ^ m[554] ^ m[556] ^ m[558] ^ m[560] ^ m[562] ^ m[564] ^ m[566] ^ m[568] ^ m[570] ^ m[572] ^ m[574] ^ m[576] ^ m[578] ^ m[580] ^ m[582] ^ m[584] ^ m[586] ^ m[588] ^ m[590] ^ m[592] ^ m[594] ^ m[596] ^ m[598] ^ m[600] ^ m[602] ^ m[604] ^ m[606] ^ m[608] ^ m[610] ^ m[612] ^ m[614] ^ m[616] ^ m[618] ^ m[620] ^ m[622] ^ m[624] ^ m[626] ^ m[628] ^ m[630] ^ m[632] ^ m[634] ^ m[636] ^ m[638] ^ m[640] ^ m[642] ^ m[644] ^ m[646] ^ m[648] ^ m[650] ^ m[652] ^ m[654] ^ m[656] ^ m[658] ^ m[660] ^ m[662] ^ m[664] ^ m[666] ^ m[668] ^ m[670] ^ m[672] ^ m[674] ^ m[676] ^ m[678] ^ m[680] ^ m[682] ^ m[684] ^ m[686] ^ m[688] ^ m[690] ^ m[692] ^ m[694] ^ m[696] ^ m[698] ^ m[700] ^ m[702] ^ m[704] ^ m[706] ^ m[708] ^ m[710] ^ m[712] ^ m[714] ^ m[716] ^ m[718] ^ m[720] ^ m[722] ^ m[724] ^ m[726] ^ m[728] ^ m[730] ^ m[732] ^ m[734] ^ m[736] ^ m[738] ^ m[740] ^ m[742] ^ m[744] ^ m[746] ^ m[748] ^ m[750] ^ m[752] ^ m[754] ^ m[756] ^ m[758] ^ m[760] ^ m[762] ^ m[764] ^ m[766] ^ m[768] ^ m[770] ^ m[772] ^ m[774] ^ m[776] ^ m[778] ^ m[780] ^ m[782] ^ m[784] ^ m[786] ^ m[788] ^ m[790] ^ m[792] ^ m[794] ^ m[796] ^ m[798] ^ m[800] ^ m[802] ^ m[804] ^ m[806] ^ m[808] ^ m[810] ^ m[812] ^ m[814] ^ m[816] ^ m[818] ^ m[820] ^ m[822] ^ m[824] ^ m[826] ^ m[828] ^ m[830] ^ m[832] ^ m[834] ^ m[836] ^ m[838] ^ m[840] ^ m[842] ^ m[844] ^ m[846] ^ m[848] ^ m[850] ^ m[852] ^ m[854] ^ m[856] ^ m[858] ^ m[860] ^ m[862] ^ m[864] ^ m[866] ^ m[868] ^ m[870] ^ m[872] ^ m[874] ^ m[876] ^ m[878] ^ m[880] ^ m[882] ^ m[884] ^ m[886] ^ m[888] ^ m[890] ^ m[892] ^ m[894] ^ m[896] ^ m[898] ^ m[900] ^ m[902] ^ m[904] ^ m[906] ^ m[908] ^ m[910] ^ m[912] ^ m[914] ^ m[916] ^ m[918] ^ m[920] ^ m[922] ^ m[924] ^ m[926] ^ m[928] ^ m[930] ^ m[932] ^ m[934] ^ m[936] ^ m[938] ^ m[940] ^ m[942] ^ m[944] ^ m[946] ^ m[948] ^ m[950] ^ m[952] ^ m[954] ^ m[956] ^ m[958] ^ m[960] ^ m[962] ^ m[964] ^ m[966] ^ m[968] ^ m[970] ^ m[972] ^ m[974] ^ m[976] ^ m[978] ^ m[980] ^ m[982] ^ m[984] ^ m[986] ^ m[988] ^ m[990] ^ m[992] ^ m[994] ^ m[996] ^ m[998] ^ m[1000] ^ m[1002] ^ m[1004] ^ m[1006] ^ m[1008] ^ m[1010] ^ m[1012] ^ m[1014] ^ m[1016] ^ m[1018] ^ m[1020] ^ m[1022] ^ m[1024] ^ m[1026] ^ m[1028] ^ m[1030] ^ m[1032] ^ m[1034] ^ m[1036] ^ m[1038] ^ m[1040] ^ m[1042] ^ m[1044] ^ m[1046] ^ m[1048] ^ m[1050] ^ m[1052] ^ m[1054] ^ m[1056] ^ m[1058] ^ m[1060] ^ m[1062] ^ m[1064] ^ m[1066] ^ m[1068] ^ m[1070] ^ m[1072] ^ m[1074] ^ m[1076] ^ m[1078] ^ m[1080] ^ m[1082] ^ m[1084] ^ m[1086] ^ m[1088] ^ m[1090] ^ m[1092] ^ m[1094] ^ m[1096] ^ m[1098] ^ m[1101] ^ m[1103] ^ m[1105] ^ m[1107] ^ m[1109] ^ m[1111] ^ m[1113] ^ m[1115] ^ m[1117] ^ m[1119] ^ m[1121] ^ m[1123] ^ m[1125] ^ m[1127] ^ m[1129] ^ m[1131] ^ m[1133] ^ m[1135] ^ m[1137] ^ m[1139] ^ m[1141] ^ m[1143] ^ m[1145] ^ m[1147] ^ m[1149] ^ m[1151] ^ m[1153] ^ m[1155] ^ m[1157] ^ m[1159] ^ m[1161] ^ m[1163] ^ m[1165] ^ m[1167] ^ m[1169] ^ m[1171] ^ m[1173] ^ m[1175] ^ m[1177] ^ m[1179] ^ m[1181] ^ m[1183] ^ m[1185] ^ m[1187] ^ m[1189] ^ m[1191] ^ m[1193] ^ m[1195] ^ m[1197] ^ m[1199] ^ m[1201] ^ m[1203] ^ m[1205] ^ m[1207] ^ m[1209] ^ m[1211] ^ m[1213] ^ m[1215] ^ m[1217] ^ m[1219] ^ m[1221] ^ m[1223] ^ m[1225] ^ m[1227] ^ m[1229] ^ m[1231] ^ m[1233] ^ m[1235] ^ m[1237] ^ m[1239] ^ m[1241] ^ m[1243] ^ m[1245] ^ m[1247] ^ m[1249] ^ m[1251] ^ m[1253] ^ m[1255] ^ m[1257] ^ m[1259] ^ m[1261] ^ m[1263] ^ m[1265] ^ m[1267] ^ m[1269] ^ m[1271] ^ m[1273] ^ m[1275] ^ m[1277] ^ m[1279] ^ m[1281] ^ m[1283] ^ m[1285] ^ m[1287] ^ m[1289] ^ m[1291] ^ m[1293] ^ m[1295] ^ m[1297] ^ m[1299] ^ m[1301] ^ m[1303] ^ m[1305] ^ m[1307] ^ m[1309] ^ m[1311] ^ m[1313] ^ m[1315] ^ m[1317] ^ m[1319] ^ m[1321] ^ m[1323] ^ m[1325] ^ m[1327] ^ m[1329] ^ m[1331] ^ m[1333] ^ m[1335] ^ m[1337] ^ m[1339] ^ m[1341] ^ m[1343] ^ m[1345] ^ m[1347] ^ m[1349] ^ m[1351] ^ m[1353] ^ m[1355] ^ m[1357] ^ m[1359] ^ m[1361] ^ m[1363] ^ m[1365] ^ m[1367] ^ m[1369] ^ m[1371] ^ m[1373] ^ m[1375] ^ m[1377] ^ m[1379] ^ m[1381] ^ m[1383] ^ m[1385] ^ m[1387] ^ m[1389] ^ m[1391] ^ m[1393] ^ m[1395] ^ m[1397] ^ m[1399] ^ m[1401] ^ m[1403] ^ m[1405] ^ m[1407] ^ m[1409] ^ m[1411] ^ m[1413] ^ m[1415] ^ m[1417] ^ m[1419] ^ m[1421] ^ m[1423] ^ m[1425] ^ m[1427] ^ m[1429] ^ m[1431] ^ m[1433] ^ m[1435] ^ m[1437] ^ m[1439] ^ m[1441] ^ m[1443] ^ m[1445] ^ m[1447] ^ m[1449] ^ m[1451] ^ m[1453] ^ m[1455] ^ m[1457] ^ m[1459] ^ m[1461] ^ m[1463] ^ m[1465] ^ m[1467] ^ m[1469] ^ m[1471] ^ m[1473] ^ m[1475] ^ m[1477] ^ m[1479] ^ m[1481] ^ m[1483] ^ m[1485] ^ m[1487] ^ m[1489] ^ m[1491] ^ m[1493] ^ m[1495] ^ m[1497] ^ m[1499] ^ m[1501] ^ m[1503] ^ m[1505] ^ m[1507] ^ m[1509] ^ m[1511] ^ m[1513] ^ m[1515] ^ m[1517] ^ m[1519] ^ m[1521] ^ m[1523] ^ m[1525] ^ m[1527] ^ m[1529] ^ m[1531] ^ m[1533] ^ m[1535] ^ m[1537] ^ m[1539] ^ m[1541] ^ m[1543] ^ m[1545] ^ m[1547] ^ m[1549] ^ m[1551] ^ m[1553] ^ m[1555] ^ m[1557] ^ m[1559] ^ m[1561] ^ m[1563] ^ m[1565] ^ m[1567] ^ m[1569] ^ m[1571] ^ m[1573] ^ m[1575] ^ m[1577] ^ m[1579] ^ m[1581] ^ m[1583] ^ m[1585] ^ m[1587] ^ m[1589] ^ m[1591] ^ m[1593] ^ m[1595] ^ m[1597] ^ m[1599] ^ m[1601] ^ m[1603] ^ m[1605] ^ m[1607] ^ m[1609] ^ m[1611] ^ m[1613] ^ m[1615] ^ m[1617] ^ m[1619] ^ m[1621] ^ m[1623] ^ m[1625] ^ m[1627] ^ m[1629] ^ m[1631] ^ m[1633] ^ m[1635] ^ m[1637] ^ m[1639] ^ m[1641] ^ m[1643] ^ m[1645] ^ m[1647] ^ m[1649] ^ m[1651] ^ m[1653] ^ m[1655] ^ m[1657] ^ m[1659] ^ m[1661] ^ m[1663] ^ m[1665] ^ m[1667] ^ m[1669] ^ m[1671] ^ m[1673] ^ m[1675] ^ m[1677] ^ m[1679] ^ m[1681] ^ m[1683] ^ m[1685] ^ m[1687] ^ m[1689] ^ m[1691] ^ m[1693] ^ m[1695] ^ m[1697] ^ m[1699] ^ m[1701] ^ m[1703] ^ m[1705] ^ m[1707] ^ m[1709] ^ m[1711] ^ m[1713] ^ m[1715] ^ m[1717] ^ m[1719] ^ m[1721] ^ m[1723] ^ m[1725] ^ m[1727] ^ m[1729] ^ m[1731] ^ m[1733] ^ m[1735] ^ m[1737] ^ m[1739] ^ m[1741] ^ m[1743] ^ m[1745] ^ m[1747] ^ m[1749] ^ m[1751] ^ m[1753] ^ m[1755] ^ m[1757] ^ m[1759] ^ m[1761] ^ m[1763] ^ m[1765] ^ m[1767] ^ m[1769] ^ m[1771] ^ m[1773] ^ m[1775] ^ m[1777] ^ m[1779] ^ m[1781] ^ m[1783] ^ m[1785] ^ m[1787] ^ m[1789] ^ m[1791] ^ m[1793] ^ m[1795] ^ m[1797] ^ m[1799] ^ m[1801] ^ m[1803] ^ m[1805] ^ m[1807] ^ m[1809] ^ m[1811] ^ m[1813] ^ m[1815] ^ m[1817] ^ m[1819] ^ m[1821] ^ m[1823] ^ m[1825] ^ m[1827] ^ m[1829] ^ m[1831] ^ m[1833] ^ m[1835] ^ m[1837] ^ m[1839] ^ m[1841] ^ m[1843] ^ m[1845] ^ m[1847] ^ m[1849] ^ m[1851] ^ m[1853] ^ m[1855] ^ m[1857] ^ m[1859] ^ m[1861] ^ m[1863] ^ m[1865] ^ m[1867] ^ m[1869] ^ m[1871] ^ m[1873] ^ m[1875] ^ m[1877] ^ m[1879] ^ m[1881] ^ m[1883] ^ m[1885] ^ m[1887] ^ m[1889] ^ m[1891] ^ m[1893] ^ m[1895] ^ m[1897] ^ m[1899] ^ m[1901] ^ m[1903] ^ m[1905] ^ m[1907] ^ m[1909] ^ m[1911] ^ m[1913] ^ m[1915] ^ m[1917] ^ m[1919] ^ m[1921] ^ m[1923] ^ m[1925] ^ m[1927] ^ m[1929] ^ m[1931] ^ m[1933] ^ m[1935] ^ m[1937] ^ m[1939] ^ m[1941] ^ m[1943] ^ m[1945] ^ m[1947] ^ m[1949] ^ m[1951] ^ m[1953] ^ m[1955] ^ m[1957] ^ m[1959] ^ m[1961] ^ m[1963] ^ m[1965] ^ m[1967] ^ m[1969] ^ m[1971] ^ m[1973] ^ m[1975] ^ m[1977] ^ m[1979] ^ m[1981] ^ m[1983] ^ m[1985] ^ m[1987] ^ m[1989] ^ m[1991] ^ m[1993] ^ m[1995] ^ m[1997] ^ m[1999] ^ m[2001] ^ m[2003] ^ m[2005] ^ m[2007] ^ m[2009] ^ m[2011] ^ m[2013] ^ m[2015] ^ m[2017] ^ m[2019] ^ m[2021] ^ m[2023] ^ m[2024] ^ m[2025] ^ m[2026] ^ m[2027] ^ m[2028] ^ m[2029] ^ m[2030] ^ m[2031] ^ m[2032] ^ m[2033] ^ m[2034];
  end else begin : gen_default_parity
    `BR_ASSERT_STATIC(invalid_parity_width_a, 1'b0)
  end

  // ri lint_check_on EXPR_ID_LIMIT

  //------
  // Concatenate message and parity bits to form the codeword.
  //------
  logic [CodewordWidth-1:0] internal_codeword;
  assign internal_codeword = {parity, m};

  //------
  // Optionally register the output signals.
  //------
  br_delay_valid #(
      .Width(CodewordWidth),
      .NumStages(RegisterOutputs == 1 ? 1 : 0),
      .EnableAssertFinalNotValid(EnableAssertFinalNotValid)
  ) br_delay_valid_outputs (
      .clk,
      .rst,
      .in_valid(data_valid_d),
      .in({internal_codeword}),
      .out_valid(enc_valid),
      .out(enc_codeword),
      .out_valid_stages(),  // unused
      .out_stages()  // unused
  );

  //------
  // Drop pad bits
  //------
  assign `BR_TRUNCATE_FROM_LSB(enc_data, enc_codeword)
  assign `BR_TRUNCATE_FROM_MSB(enc_parity, enc_codeword)
  if (OutputWidth < CodewordWidth) begin : gen_unused_out
    `BR_UNUSED_NAMED(unused_out, enc_codeword[MessageWidth-1 : DataWidth])
  end

  //------------------------------------------
  // Implementation checks
  //------------------------------------------
  `BR_ASSERT_IMPL(latency_a, data_valid |-> ##Latency enc_valid)

  // verilog_lint: waive-stop line-length
  // verilog_format: on

endmodule : br_ecc_secded_encoder
