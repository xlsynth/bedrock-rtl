// Copyright 2024 The Bedrock-RTL Authors
//
// Licensed under the Apache License, Version 2.0 (the "License");
// Copyright 2024 The Bedrock-RTL Authors
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//     http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.


// verilog_format: off
// verilog_lint: waive-start line-length

// Bedrock-RTL Single-Error-Correcting, Double-Error-Detecting (SECDED - Hsiao) Encoder
//
// Encodes a message using a single-error-correcting, double-error-detecting
// linear block code in systematic form (in layperson's terms: a Hsiao SECDED [1] encoder,
// closely related to Hamming codes).
//
// Systematic form means that the codeword is formed by appending the
// calculated parity bits to the message, i.e., the code has the property
// that the message bits are 1:1 with a slice of bits in the codeword (if they
// have not been corrupted).
//
// In Bedrock ECC libs, our convention is to always append the parity bits on
// the MSbs:
//     codeword == {parity, message}
//
// This module has parameterizable latency. By default, it is purely combinational,
// but it can have up to 2 cycles of delay (RegisterInputs and RegisterOutputs).
// The initiation interval is always 1 cycle.
//
// Any data width >= 1 is supported. It is internally zero-padded up to
// the nearest power-of-2 message width before being encoded. The following
// table outlines the number of parity bits required for different message widths.
//
// | Message Width (k) | Parity Width (r) | Codeword Width (n)|
// |-------------------|------------------|-------------------|
// | 4                 | 4                | 8                 |
// | 8                 | 5                | 13                |
// | 16                | 6                | 22                |
// | 32                | 7                | 39                |
// | 64                | 8                | 72                |
// | 128               | 9                | 137               |
// | 256               | 10               | 266               |
// | 512               | 11               | 523               |
// | 1024              | 12               | 1036              |
//
// The number of parity bits must be one of the values in the table above
// or the module will not elaborate.
//
// References:
// [1] https://ieeexplore.ieee.org/abstract/document/5391627

`include "br_asserts.svh"
`include "br_asserts_internal.svh"

module br_ecc_secded_encoder #(
    parameter int DataWidth = 1,  // Must be at least 1
    parameter int ParityWidth = 4,  // Must be at least 4 and at most 12
    // If 1, then insert a pipeline register at the input.
    parameter bit RegisterInputs = 0,
    // If 1, then insert a pipeline register at the output.
    parameter bit RegisterOutputs = 0,
    localparam int MessageWidth = 2 ** $clog2(DataWidth),
    localparam int CodewordWidth = MessageWidth + ParityWidth
) (
    // Positive edge-triggered clock.
    input  logic                     clk,
    // Synchronous active-high reset.
    input  logic                     rst,
    input  logic                     data_valid,
    input  logic [    DataWidth-1:0] data,
    output logic                     enc_valid,
    output logic [CodewordWidth-1:0] enc_codeword
);

  // ri lint_check_waive PARAM_NOT_USED
  localparam int Latency = RegisterOutputs ? 1 : 0;

  //------------------------------------------
  // Integration checks
  //------------------------------------------
  `BR_ASSERT_STATIC(message_width_gte_1_a, DataWidth >= 1)
  `BR_ASSERT_STATIC(parity_width_gte_4_a, ParityWidth >= 4)
  `BR_ASSERT_STATIC(parity_width_lte_12_a, ParityWidth <= 12)
  `BR_ASSERT_STATIC(message_width_is_power_of_2_a, br_math::is_power_of_2(MessageWidth))

  //------------------------------------------
  // Implementation
  //------------------------------------------

  //------
  // Optionally register the input signals.
  //------
  logic data_valid_d;
  logic [DataWidth-1:0] data_d;

  br_delay_valid #(
      .Width(DataWidth),
      .NumStages(RegisterInputs == 1 ? 1 : 0)
  ) br_delay_valid_inputs (
      .clk,
      .rst,
      .in_valid(data_valid),
      .in(data),
      .out_valid(data_valid_d),
      .out(data_d),
      .out_valid_stages(),  // unused
      .out_stages()  // unused
  );

  //------
  // Pad the data to the nearest power of 2 message width.
  //------

  localparam int PadWidth = MessageWidth - DataWidth;
  logic [MessageWidth-1:0] m;

  if (PadWidth > 0) begin : gen_pad
    assign m = { {PadWidth{1'b0} }, data_d};
  end else begin : gen_no_pad
    assign m = data_d;
  end

  //------
  // Compute parity bits.
  //------
  logic [ParityWidth-1:0] parity;

  // ri lint_check_off EXPR_ID_LIMIT

  if ((CodewordWidth == 4) && (MessageWidth == 4)) begin : gen_8_4
    `BR_ASSERT_STATIC(parity_width_matches_a, ParityWidth == 4)
    assign parity[0] = m[1] ^ m[2] ^ m[3];
    assign parity[1] = m[0] ^ m[2] ^ m[3];
    assign parity[2] = m[0] ^ m[1] ^ m[3];
    assign parity[3] = m[0] ^ m[1] ^ m[2];
  end else if ((CodewordWidth == 13) && (MessageWidth == 8)) begin : gen_13_8
    `BR_ASSERT_STATIC(parity_width_matches_a, ParityWidth == 5)
    assign parity[0] = m[4] ^ m[5] ^ m[6] ^ m[7];
    assign parity[1] = m[1] ^ m[2] ^ m[3] ^ m[7];
    assign parity[2] = m[0] ^ m[2] ^ m[3] ^ m[5] ^ m[6];
    assign parity[3] = m[0] ^ m[1] ^ m[3] ^ m[4] ^ m[6];
    assign parity[4] = m[0] ^ m[1] ^ m[2] ^ m[4] ^ m[5] ^ m[7];
  end else if ((CodewordWidth == 22) && (MessageWidth == 16)) begin : gen_22_16
    `BR_ASSERT_STATIC(parity_width_matches_a, ParityWidth == 6)
    assign parity[0] = m[10] ^ m[11] ^ m[12] ^ m[13] ^ m[14] ^ m[15];
    assign parity[1] = m[4] ^ m[5] ^ m[6] ^ m[7] ^ m[8] ^ m[9];
    assign parity[2] = m[1] ^ m[2] ^ m[3] ^ m[7] ^ m[8] ^ m[9] ^ m[13] ^ m[14] ^ m[15];
    assign parity[3] = m[0] ^ m[2] ^ m[3] ^ m[5] ^ m[6] ^ m[9] ^ m[11] ^ m[12] ^ m[15];
    assign parity[4] = m[0] ^ m[1] ^ m[3] ^ m[4] ^ m[6] ^ m[8] ^ m[10] ^ m[12] ^ m[14];
    assign parity[5] = m[0] ^ m[1] ^ m[2] ^ m[4] ^ m[5] ^ m[7] ^ m[10] ^ m[11] ^ m[13];
  end else if ((CodewordWidth == 39) && (MessageWidth == 32)) begin : gen_39_32
    `BR_ASSERT_STATIC(parity_width_matches_a, ParityWidth == 7)
    assign parity[0] = m[20] ^ m[21] ^ m[22] ^ m[23] ^ m[24] ^ m[25] ^ m[26] ^ m[27] ^ m[28] ^ m[29] ^ m[30] ^ m[31];
    assign parity[1] = m[10] ^ m[11] ^ m[12] ^ m[13] ^ m[14] ^ m[15] ^ m[16] ^ m[17] ^ m[18] ^ m[19] ^ m[30] ^ m[31];
    assign parity[2] = m[4] ^ m[5] ^ m[6] ^ m[7] ^ m[8] ^ m[9] ^ m[16] ^ m[17] ^ m[18] ^ m[19] ^ m[26] ^ m[27] ^ m[28] ^ m[29];
    assign parity[3] = m[1] ^ m[2] ^ m[3] ^ m[7] ^ m[8] ^ m[9] ^ m[13] ^ m[14] ^ m[15] ^ m[19] ^ m[23] ^ m[24] ^ m[25] ^ m[29];
    assign parity[4] = m[0] ^ m[2] ^ m[3] ^ m[5] ^ m[6] ^ m[9] ^ m[11] ^ m[12] ^ m[15] ^ m[18] ^ m[21] ^ m[22] ^ m[25] ^ m[28];
    assign parity[5] = m[0] ^ m[1] ^ m[3] ^ m[4] ^ m[6] ^ m[8] ^ m[10] ^ m[12] ^ m[14] ^ m[17] ^ m[20] ^ m[22] ^ m[24] ^ m[27] ^ m[31];
    assign parity[6] = m[0] ^ m[1] ^ m[2] ^ m[4] ^ m[5] ^ m[7] ^ m[10] ^ m[11] ^ m[13] ^ m[16] ^ m[20] ^ m[21] ^ m[23] ^ m[26] ^ m[30];
  end else if ((CodewordWidth == 72) && (MessageWidth == 64)) begin : gen_72_64
    `BR_ASSERT_STATIC(parity_width_matches_a, ParityWidth == 8)
    assign parity[0] = m[35] ^ m[36] ^ m[37] ^ m[38] ^ m[39] ^ m[40] ^ m[41] ^ m[42] ^ m[43] ^ m[44] ^ m[45] ^ m[46] ^ m[47] ^ m[48] ^ m[49] ^ m[50] ^ m[51] ^ m[52] ^ m[53] ^ m[54] ^ m[55];
    assign parity[1] = m[20] ^ m[21] ^ m[22] ^ m[23] ^ m[24] ^ m[25] ^ m[26] ^ m[27] ^ m[28] ^ m[29] ^ m[30] ^ m[31] ^ m[32] ^ m[33] ^ m[34] ^ m[50] ^ m[51] ^ m[52] ^ m[53] ^ m[54] ^ m[55] ^ m[62] ^ m[63];
    assign parity[2] = m[10] ^ m[11] ^ m[12] ^ m[13] ^ m[14] ^ m[15] ^ m[16] ^ m[17] ^ m[18] ^ m[19] ^ m[30] ^ m[31] ^ m[32] ^ m[33] ^ m[34] ^ m[45] ^ m[46] ^ m[47] ^ m[48] ^ m[49] ^ m[55] ^ m[57] ^ m[58] ^ m[59] ^ m[60] ^ m[61];
    assign parity[3] = m[4] ^ m[5] ^ m[6] ^ m[7] ^ m[8] ^ m[9] ^ m[16] ^ m[17] ^ m[18] ^ m[19] ^ m[26] ^ m[27] ^ m[28] ^ m[29] ^ m[34] ^ m[41] ^ m[42] ^ m[43] ^ m[44] ^ m[49] ^ m[54] ^ m[56] ^ m[58] ^ m[59] ^ m[60] ^ m[61] ^ m[63];
    assign parity[4] = m[1] ^ m[2] ^ m[3] ^ m[7] ^ m[8] ^ m[9] ^ m[13] ^ m[14] ^ m[15] ^ m[19] ^ m[23] ^ m[24] ^ m[25] ^ m[29] ^ m[33] ^ m[38] ^ m[39] ^ m[40] ^ m[44] ^ m[48] ^ m[53] ^ m[56] ^ m[57] ^ m[59] ^ m[60] ^ m[61] ^ m[62];
    assign parity[5] = m[0] ^ m[2] ^ m[3] ^ m[5] ^ m[6] ^ m[9] ^ m[11] ^ m[12] ^ m[15] ^ m[18] ^ m[21] ^ m[22] ^ m[25] ^ m[28] ^ m[32] ^ m[36] ^ m[37] ^ m[40] ^ m[43] ^ m[47] ^ m[52] ^ m[56] ^ m[57] ^ m[58] ^ m[60] ^ m[61] ^ m[62] ^ m[63];
    assign parity[6] = m[0] ^ m[1] ^ m[3] ^ m[4] ^ m[6] ^ m[8] ^ m[10] ^ m[12] ^ m[14] ^ m[17] ^ m[20] ^ m[22] ^ m[24] ^ m[27] ^ m[31] ^ m[35] ^ m[37] ^ m[39] ^ m[42] ^ m[46] ^ m[51] ^ m[56] ^ m[57] ^ m[58] ^ m[59] ^ m[61] ^ m[62] ^ m[63];
    assign parity[7] = m[0] ^ m[1] ^ m[2] ^ m[4] ^ m[5] ^ m[7] ^ m[10] ^ m[11] ^ m[13] ^ m[16] ^ m[20] ^ m[21] ^ m[23] ^ m[26] ^ m[30] ^ m[35] ^ m[36] ^ m[38] ^ m[41] ^ m[45] ^ m[50] ^ m[56] ^ m[57] ^ m[58] ^ m[59] ^ m[60] ^ m[62] ^ m[63];
  end else if ((CodewordWidth == 137) && (MessageWidth == 128)) begin : gen_137_128
    `BR_ASSERT_STATIC(parity_width_matches_a, ParityWidth == 9)
    assign parity[0] = m[56] ^ m[57] ^ m[58] ^ m[59] ^ m[60] ^ m[61] ^ m[62] ^ m[63] ^ m[64] ^ m[65] ^ m[66] ^ m[67] ^ m[68] ^ m[69] ^ m[70] ^ m[71] ^ m[72] ^ m[73] ^ m[74] ^ m[75] ^ m[76] ^ m[77] ^ m[78] ^ m[79] ^ m[80] ^ m[81] ^ m[82] ^ m[83];
    assign parity[1] = m[35] ^ m[36] ^ m[37] ^ m[38] ^ m[39] ^ m[40] ^ m[41] ^ m[42] ^ m[43] ^ m[44] ^ m[45] ^ m[46] ^ m[47] ^ m[48] ^ m[49] ^ m[50] ^ m[51] ^ m[52] ^ m[53] ^ m[54] ^ m[55] ^ m[77] ^ m[78] ^ m[79] ^ m[80] ^ m[81] ^ m[82] ^ m[83] ^ m[105] ^ m[106] ^ m[107] ^ m[108] ^ m[109] ^ m[110] ^ m[111] ^ m[112] ^ m[113] ^ m[114] ^ m[115] ^ m[116] ^ m[117] ^ m[118] ^ m[119] ^ m[120] ^ m[121] ^ m[122] ^ m[123] ^ m[124] ^ m[125] ^ m[126] ^ m[127];
    assign parity[2] = m[20] ^ m[21] ^ m[22] ^ m[23] ^ m[24] ^ m[25] ^ m[26] ^ m[27] ^ m[28] ^ m[29] ^ m[30] ^ m[31] ^ m[32] ^ m[33] ^ m[34] ^ m[50] ^ m[51] ^ m[52] ^ m[53] ^ m[54] ^ m[55] ^ m[71] ^ m[72] ^ m[73] ^ m[74] ^ m[75] ^ m[76] ^ m[83] ^ m[90] ^ m[91] ^ m[92] ^ m[93] ^ m[94] ^ m[95] ^ m[96] ^ m[97] ^ m[98] ^ m[99] ^ m[100] ^ m[101] ^ m[102] ^ m[103] ^ m[104] ^ m[120] ^ m[121] ^ m[122] ^ m[123] ^ m[124] ^ m[125] ^ m[126] ^ m[127];
    assign parity[3] = m[10] ^ m[11] ^ m[12] ^ m[13] ^ m[14] ^ m[15] ^ m[16] ^ m[17] ^ m[18] ^ m[19] ^ m[30] ^ m[31] ^ m[32] ^ m[33] ^ m[34] ^ m[45] ^ m[46] ^ m[47] ^ m[48] ^ m[49] ^ m[55] ^ m[66] ^ m[67] ^ m[68] ^ m[69] ^ m[70] ^ m[76] ^ m[82] ^ m[85] ^ m[86] ^ m[87] ^ m[88] ^ m[89] ^ m[95] ^ m[96] ^ m[97] ^ m[98] ^ m[99] ^ m[100] ^ m[101] ^ m[102] ^ m[103] ^ m[104] ^ m[110] ^ m[111] ^ m[112] ^ m[113] ^ m[114] ^ m[115] ^ m[116] ^ m[117] ^ m[118] ^ m[119];
    assign parity[4] = m[4] ^ m[5] ^ m[6] ^ m[7] ^ m[8] ^ m[9] ^ m[16] ^ m[17] ^ m[18] ^ m[19] ^ m[26] ^ m[27] ^ m[28] ^ m[29] ^ m[34] ^ m[41] ^ m[42] ^ m[43] ^ m[44] ^ m[49] ^ m[54] ^ m[62] ^ m[63] ^ m[64] ^ m[65] ^ m[70] ^ m[75] ^ m[81] ^ m[84] ^ m[86] ^ m[87] ^ m[88] ^ m[89] ^ m[91] ^ m[92] ^ m[93] ^ m[94] ^ m[99] ^ m[100] ^ m[101] ^ m[102] ^ m[103] ^ m[104] ^ m[106] ^ m[107] ^ m[108] ^ m[109] ^ m[114] ^ m[115] ^ m[116] ^ m[117] ^ m[118] ^ m[119] ^ m[124] ^ m[125] ^ m[126] ^ m[127];
    assign parity[5] = m[1] ^ m[2] ^ m[3] ^ m[7] ^ m[8] ^ m[9] ^ m[13] ^ m[14] ^ m[15] ^ m[19] ^ m[23] ^ m[24] ^ m[25] ^ m[29] ^ m[33] ^ m[38] ^ m[39] ^ m[40] ^ m[44] ^ m[48] ^ m[53] ^ m[59] ^ m[60] ^ m[61] ^ m[65] ^ m[69] ^ m[74] ^ m[80] ^ m[84] ^ m[85] ^ m[87] ^ m[88] ^ m[89] ^ m[90] ^ m[92] ^ m[93] ^ m[94] ^ m[96] ^ m[97] ^ m[98] ^ m[102] ^ m[103] ^ m[104] ^ m[105] ^ m[107] ^ m[108] ^ m[109] ^ m[111] ^ m[112] ^ m[113] ^ m[117] ^ m[118] ^ m[119] ^ m[121] ^ m[122] ^ m[123] ^ m[127];
    assign parity[6] = m[0] ^ m[2] ^ m[3] ^ m[5] ^ m[6] ^ m[9] ^ m[11] ^ m[12] ^ m[15] ^ m[18] ^ m[21] ^ m[22] ^ m[25] ^ m[28] ^ m[32] ^ m[36] ^ m[37] ^ m[40] ^ m[43] ^ m[47] ^ m[52] ^ m[57] ^ m[58] ^ m[61] ^ m[64] ^ m[68] ^ m[73] ^ m[79] ^ m[84] ^ m[85] ^ m[86] ^ m[88] ^ m[89] ^ m[90] ^ m[91] ^ m[93] ^ m[94] ^ m[95] ^ m[97] ^ m[98] ^ m[100] ^ m[101] ^ m[104] ^ m[105] ^ m[106] ^ m[108] ^ m[109] ^ m[110] ^ m[112] ^ m[113] ^ m[115] ^ m[116] ^ m[119] ^ m[120] ^ m[122] ^ m[123] ^ m[125] ^ m[126];
    assign parity[7] = m[0] ^ m[1] ^ m[3] ^ m[4] ^ m[6] ^ m[8] ^ m[10] ^ m[12] ^ m[14] ^ m[17] ^ m[20] ^ m[22] ^ m[24] ^ m[27] ^ m[31] ^ m[35] ^ m[37] ^ m[39] ^ m[42] ^ m[46] ^ m[51] ^ m[56] ^ m[58] ^ m[60] ^ m[63] ^ m[67] ^ m[72] ^ m[78] ^ m[84] ^ m[85] ^ m[86] ^ m[87] ^ m[89] ^ m[90] ^ m[91] ^ m[92] ^ m[94] ^ m[95] ^ m[96] ^ m[98] ^ m[99] ^ m[101] ^ m[103] ^ m[105] ^ m[106] ^ m[107] ^ m[109] ^ m[110] ^ m[111] ^ m[113] ^ m[114] ^ m[116] ^ m[118] ^ m[120] ^ m[121] ^ m[123] ^ m[124] ^ m[126];
    assign parity[8] = m[0] ^ m[1] ^ m[2] ^ m[4] ^ m[5] ^ m[7] ^ m[10] ^ m[11] ^ m[13] ^ m[16] ^ m[20] ^ m[21] ^ m[23] ^ m[26] ^ m[30] ^ m[35] ^ m[36] ^ m[38] ^ m[41] ^ m[45] ^ m[50] ^ m[56] ^ m[57] ^ m[59] ^ m[62] ^ m[66] ^ m[71] ^ m[77] ^ m[84] ^ m[85] ^ m[86] ^ m[87] ^ m[88] ^ m[90] ^ m[91] ^ m[92] ^ m[93] ^ m[95] ^ m[96] ^ m[97] ^ m[99] ^ m[100] ^ m[102] ^ m[105] ^ m[106] ^ m[107] ^ m[108] ^ m[110] ^ m[111] ^ m[112] ^ m[114] ^ m[115] ^ m[117] ^ m[120] ^ m[121] ^ m[122] ^ m[124] ^ m[125] ^ m[127];
  end else if ((CodewordWidth == 266) && (MessageWidth == 256)) begin : gen_266_256
    `BR_ASSERT_STATIC(parity_width_matches_a, ParityWidth == 10)
    assign parity[0] = m[84] ^ m[85] ^ m[86] ^ m[87] ^ m[88] ^ m[89] ^ m[90] ^ m[91] ^ m[92] ^ m[93] ^ m[94] ^ m[95] ^ m[96] ^ m[97] ^ m[98] ^ m[99] ^ m[100] ^ m[101] ^ m[102] ^ m[103] ^ m[104] ^ m[105] ^ m[106] ^ m[107] ^ m[108] ^ m[109] ^ m[110] ^ m[111] ^ m[112] ^ m[113] ^ m[114] ^ m[115] ^ m[116] ^ m[117] ^ m[118] ^ m[119] ^ m[246] ^ m[247] ^ m[248] ^ m[249] ^ m[250] ^ m[251] ^ m[252] ^ m[253] ^ m[254] ^ m[255];
    assign parity[1] = m[56] ^ m[57] ^ m[58] ^ m[59] ^ m[60] ^ m[61] ^ m[62] ^ m[63] ^ m[64] ^ m[65] ^ m[66] ^ m[67] ^ m[68] ^ m[69] ^ m[70] ^ m[71] ^ m[72] ^ m[73] ^ m[74] ^ m[75] ^ m[76] ^ m[77] ^ m[78] ^ m[79] ^ m[80] ^ m[81] ^ m[82] ^ m[83] ^ m[112] ^ m[113] ^ m[114] ^ m[115] ^ m[116] ^ m[117] ^ m[118] ^ m[119] ^ m[176] ^ m[177] ^ m[178] ^ m[179] ^ m[180] ^ m[181] ^ m[182] ^ m[183] ^ m[184] ^ m[185] ^ m[186] ^ m[187] ^ m[188] ^ m[189] ^ m[190] ^ m[191] ^ m[192] ^ m[193] ^ m[194] ^ m[195] ^ m[196] ^ m[197] ^ m[198] ^ m[199] ^ m[200] ^ m[201] ^ m[202] ^ m[203] ^ m[204] ^ m[205] ^ m[206] ^ m[207] ^ m[208] ^ m[209] ^ m[210] ^ m[211] ^ m[212] ^ m[213] ^ m[214] ^ m[215] ^ m[216] ^ m[217] ^ m[218] ^ m[219] ^ m[220] ^ m[221] ^ m[222] ^ m[223] ^ m[224] ^ m[225] ^ m[226] ^ m[227] ^ m[228] ^ m[229] ^ m[230] ^ m[231] ^ m[232] ^ m[233] ^ m[234] ^ m[235] ^ m[236] ^ m[237] ^ m[238] ^ m[239] ^ m[240] ^ m[241] ^ m[242] ^ m[243] ^ m[244] ^ m[245];
    assign parity[2] = m[35] ^ m[36] ^ m[37] ^ m[38] ^ m[39] ^ m[40] ^ m[41] ^ m[42] ^ m[43] ^ m[44] ^ m[45] ^ m[46] ^ m[47] ^ m[48] ^ m[49] ^ m[50] ^ m[51] ^ m[52] ^ m[53] ^ m[54] ^ m[55] ^ m[77] ^ m[78] ^ m[79] ^ m[80] ^ m[81] ^ m[82] ^ m[83] ^ m[105] ^ m[106] ^ m[107] ^ m[108] ^ m[109] ^ m[110] ^ m[111] ^ m[119] ^ m[141] ^ m[142] ^ m[143] ^ m[144] ^ m[145] ^ m[146] ^ m[147] ^ m[148] ^ m[149] ^ m[150] ^ m[151] ^ m[152] ^ m[153] ^ m[154] ^ m[155] ^ m[156] ^ m[157] ^ m[158] ^ m[159] ^ m[160] ^ m[161] ^ m[162] ^ m[163] ^ m[164] ^ m[165] ^ m[166] ^ m[167] ^ m[168] ^ m[169] ^ m[170] ^ m[171] ^ m[172] ^ m[173] ^ m[174] ^ m[175] ^ m[211] ^ m[212] ^ m[213] ^ m[214] ^ m[215] ^ m[216] ^ m[217] ^ m[218] ^ m[219] ^ m[220] ^ m[221] ^ m[222] ^ m[223] ^ m[224] ^ m[225] ^ m[226] ^ m[227] ^ m[228] ^ m[229] ^ m[230] ^ m[231] ^ m[232] ^ m[233] ^ m[234] ^ m[235] ^ m[236] ^ m[237] ^ m[238] ^ m[239] ^ m[240] ^ m[241] ^ m[242] ^ m[243] ^ m[244] ^ m[245];
    assign parity[3] = m[20] ^ m[21] ^ m[22] ^ m[23] ^ m[24] ^ m[25] ^ m[26] ^ m[27] ^ m[28] ^ m[29] ^ m[30] ^ m[31] ^ m[32] ^ m[33] ^ m[34] ^ m[50] ^ m[51] ^ m[52] ^ m[53] ^ m[54] ^ m[55] ^ m[71] ^ m[72] ^ m[73] ^ m[74] ^ m[75] ^ m[76] ^ m[83] ^ m[99] ^ m[100] ^ m[101] ^ m[102] ^ m[103] ^ m[104] ^ m[111] ^ m[118] ^ m[126] ^ m[127] ^ m[128] ^ m[129] ^ m[130] ^ m[131] ^ m[132] ^ m[133] ^ m[134] ^ m[135] ^ m[136] ^ m[137] ^ m[138] ^ m[139] ^ m[140] ^ m[156] ^ m[157] ^ m[158] ^ m[159] ^ m[160] ^ m[161] ^ m[162] ^ m[163] ^ m[164] ^ m[165] ^ m[166] ^ m[167] ^ m[168] ^ m[169] ^ m[170] ^ m[171] ^ m[172] ^ m[173] ^ m[174] ^ m[175] ^ m[191] ^ m[192] ^ m[193] ^ m[194] ^ m[195] ^ m[196] ^ m[197] ^ m[198] ^ m[199] ^ m[200] ^ m[201] ^ m[202] ^ m[203] ^ m[204] ^ m[205] ^ m[206] ^ m[207] ^ m[208] ^ m[209] ^ m[210] ^ m[231] ^ m[232] ^ m[233] ^ m[234] ^ m[235] ^ m[236] ^ m[237] ^ m[238] ^ m[239] ^ m[240] ^ m[241] ^ m[242] ^ m[243] ^ m[244] ^ m[245];
    assign parity[4] = m[10] ^ m[11] ^ m[12] ^ m[13] ^ m[14] ^ m[15] ^ m[16] ^ m[17] ^ m[18] ^ m[19] ^ m[30] ^ m[31] ^ m[32] ^ m[33] ^ m[34] ^ m[45] ^ m[46] ^ m[47] ^ m[48] ^ m[49] ^ m[55] ^ m[66] ^ m[67] ^ m[68] ^ m[69] ^ m[70] ^ m[76] ^ m[82] ^ m[94] ^ m[95] ^ m[96] ^ m[97] ^ m[98] ^ m[104] ^ m[110] ^ m[117] ^ m[121] ^ m[122] ^ m[123] ^ m[124] ^ m[125] ^ m[131] ^ m[132] ^ m[133] ^ m[134] ^ m[135] ^ m[136] ^ m[137] ^ m[138] ^ m[139] ^ m[140] ^ m[146] ^ m[147] ^ m[148] ^ m[149] ^ m[150] ^ m[151] ^ m[152] ^ m[153] ^ m[154] ^ m[155] ^ m[166] ^ m[167] ^ m[168] ^ m[169] ^ m[170] ^ m[171] ^ m[172] ^ m[173] ^ m[174] ^ m[175] ^ m[181] ^ m[182] ^ m[183] ^ m[184] ^ m[185] ^ m[186] ^ m[187] ^ m[188] ^ m[189] ^ m[190] ^ m[201] ^ m[202] ^ m[203] ^ m[204] ^ m[205] ^ m[206] ^ m[207] ^ m[208] ^ m[209] ^ m[210] ^ m[221] ^ m[222] ^ m[223] ^ m[224] ^ m[225] ^ m[226] ^ m[227] ^ m[228] ^ m[229] ^ m[230] ^ m[241] ^ m[242] ^ m[243] ^ m[244] ^ m[245] ^ m[251] ^ m[252] ^ m[253] ^ m[254] ^ m[255];
    assign parity[5] = m[4] ^ m[5] ^ m[6] ^ m[7] ^ m[8] ^ m[9] ^ m[16] ^ m[17] ^ m[18] ^ m[19] ^ m[26] ^ m[27] ^ m[28] ^ m[29] ^ m[34] ^ m[41] ^ m[42] ^ m[43] ^ m[44] ^ m[49] ^ m[54] ^ m[62] ^ m[63] ^ m[64] ^ m[65] ^ m[70] ^ m[75] ^ m[81] ^ m[90] ^ m[91] ^ m[92] ^ m[93] ^ m[98] ^ m[103] ^ m[109] ^ m[116] ^ m[120] ^ m[122] ^ m[123] ^ m[124] ^ m[125] ^ m[127] ^ m[128] ^ m[129] ^ m[130] ^ m[135] ^ m[136] ^ m[137] ^ m[138] ^ m[139] ^ m[140] ^ m[142] ^ m[143] ^ m[144] ^ m[145] ^ m[150] ^ m[151] ^ m[152] ^ m[153] ^ m[154] ^ m[155] ^ m[160] ^ m[161] ^ m[162] ^ m[163] ^ m[164] ^ m[165] ^ m[172] ^ m[173] ^ m[174] ^ m[175] ^ m[177] ^ m[178] ^ m[179] ^ m[180] ^ m[185] ^ m[186] ^ m[187] ^ m[188] ^ m[189] ^ m[190] ^ m[195] ^ m[196] ^ m[197] ^ m[198] ^ m[199] ^ m[200] ^ m[207] ^ m[208] ^ m[209] ^ m[210] ^ m[215] ^ m[216] ^ m[217] ^ m[218] ^ m[219] ^ m[220] ^ m[227] ^ m[228] ^ m[229] ^ m[230] ^ m[237] ^ m[238] ^ m[239] ^ m[240] ^ m[245] ^ m[247] ^ m[248] ^ m[249] ^ m[250] ^ m[255];
    assign parity[6] = m[1] ^ m[2] ^ m[3] ^ m[7] ^ m[8] ^ m[9] ^ m[13] ^ m[14] ^ m[15] ^ m[19] ^ m[23] ^ m[24] ^ m[25] ^ m[29] ^ m[33] ^ m[38] ^ m[39] ^ m[40] ^ m[44] ^ m[48] ^ m[53] ^ m[59] ^ m[60] ^ m[61] ^ m[65] ^ m[69] ^ m[74] ^ m[80] ^ m[87] ^ m[88] ^ m[89] ^ m[93] ^ m[97] ^ m[102] ^ m[108] ^ m[115] ^ m[120] ^ m[121] ^ m[123] ^ m[124] ^ m[125] ^ m[126] ^ m[128] ^ m[129] ^ m[130] ^ m[132] ^ m[133] ^ m[134] ^ m[138] ^ m[139] ^ m[140] ^ m[141] ^ m[143] ^ m[144] ^ m[145] ^ m[147] ^ m[148] ^ m[149] ^ m[153] ^ m[154] ^ m[155] ^ m[157] ^ m[158] ^ m[159] ^ m[163] ^ m[164] ^ m[165] ^ m[169] ^ m[170] ^ m[171] ^ m[175] ^ m[176] ^ m[178] ^ m[179] ^ m[180] ^ m[182] ^ m[183] ^ m[184] ^ m[188] ^ m[189] ^ m[190] ^ m[192] ^ m[193] ^ m[194] ^ m[198] ^ m[199] ^ m[200] ^ m[204] ^ m[205] ^ m[206] ^ m[210] ^ m[212] ^ m[213] ^ m[214] ^ m[218] ^ m[219] ^ m[220] ^ m[224] ^ m[225] ^ m[226] ^ m[230] ^ m[234] ^ m[235] ^ m[236] ^ m[240] ^ m[244] ^ m[246] ^ m[248] ^ m[249] ^ m[250] ^ m[252] ^ m[253] ^ m[254];
    assign parity[7] = m[0] ^ m[2] ^ m[3] ^ m[5] ^ m[6] ^ m[9] ^ m[11] ^ m[12] ^ m[15] ^ m[18] ^ m[21] ^ m[22] ^ m[25] ^ m[28] ^ m[32] ^ m[36] ^ m[37] ^ m[40] ^ m[43] ^ m[47] ^ m[52] ^ m[57] ^ m[58] ^ m[61] ^ m[64] ^ m[68] ^ m[73] ^ m[79] ^ m[85] ^ m[86] ^ m[89] ^ m[92] ^ m[96] ^ m[101] ^ m[107] ^ m[114] ^ m[120] ^ m[121] ^ m[122] ^ m[124] ^ m[125] ^ m[126] ^ m[127] ^ m[129] ^ m[130] ^ m[131] ^ m[133] ^ m[134] ^ m[136] ^ m[137] ^ m[140] ^ m[141] ^ m[142] ^ m[144] ^ m[145] ^ m[146] ^ m[148] ^ m[149] ^ m[151] ^ m[152] ^ m[155] ^ m[156] ^ m[158] ^ m[159] ^ m[161] ^ m[162] ^ m[165] ^ m[167] ^ m[168] ^ m[171] ^ m[174] ^ m[176] ^ m[177] ^ m[179] ^ m[180] ^ m[181] ^ m[183] ^ m[184] ^ m[186] ^ m[187] ^ m[190] ^ m[191] ^ m[193] ^ m[194] ^ m[196] ^ m[197] ^ m[200] ^ m[202] ^ m[203] ^ m[206] ^ m[209] ^ m[211] ^ m[213] ^ m[214] ^ m[216] ^ m[217] ^ m[220] ^ m[222] ^ m[223] ^ m[226] ^ m[229] ^ m[232] ^ m[233] ^ m[236] ^ m[239] ^ m[243] ^ m[246] ^ m[247] ^ m[249] ^ m[250] ^ m[251] ^ m[253] ^ m[254];
    assign parity[8] = m[0] ^ m[1] ^ m[3] ^ m[4] ^ m[6] ^ m[8] ^ m[10] ^ m[12] ^ m[14] ^ m[17] ^ m[20] ^ m[22] ^ m[24] ^ m[27] ^ m[31] ^ m[35] ^ m[37] ^ m[39] ^ m[42] ^ m[46] ^ m[51] ^ m[56] ^ m[58] ^ m[60] ^ m[63] ^ m[67] ^ m[72] ^ m[78] ^ m[84] ^ m[86] ^ m[88] ^ m[91] ^ m[95] ^ m[100] ^ m[106] ^ m[113] ^ m[120] ^ m[121] ^ m[122] ^ m[123] ^ m[125] ^ m[126] ^ m[127] ^ m[128] ^ m[130] ^ m[131] ^ m[132] ^ m[134] ^ m[135] ^ m[137] ^ m[139] ^ m[141] ^ m[142] ^ m[143] ^ m[145] ^ m[146] ^ m[147] ^ m[149] ^ m[150] ^ m[152] ^ m[154] ^ m[156] ^ m[157] ^ m[159] ^ m[160] ^ m[162] ^ m[164] ^ m[166] ^ m[168] ^ m[170] ^ m[173] ^ m[176] ^ m[177] ^ m[178] ^ m[180] ^ m[181] ^ m[182] ^ m[184] ^ m[185] ^ m[187] ^ m[189] ^ m[191] ^ m[192] ^ m[194] ^ m[195] ^ m[197] ^ m[199] ^ m[201] ^ m[203] ^ m[205] ^ m[208] ^ m[211] ^ m[212] ^ m[214] ^ m[215] ^ m[217] ^ m[219] ^ m[221] ^ m[223] ^ m[225] ^ m[228] ^ m[231] ^ m[233] ^ m[235] ^ m[238] ^ m[242] ^ m[246] ^ m[247] ^ m[248] ^ m[250] ^ m[251] ^ m[252] ^ m[254] ^ m[255];
    assign parity[9] = m[0] ^ m[1] ^ m[2] ^ m[4] ^ m[5] ^ m[7] ^ m[10] ^ m[11] ^ m[13] ^ m[16] ^ m[20] ^ m[21] ^ m[23] ^ m[26] ^ m[30] ^ m[35] ^ m[36] ^ m[38] ^ m[41] ^ m[45] ^ m[50] ^ m[56] ^ m[57] ^ m[59] ^ m[62] ^ m[66] ^ m[71] ^ m[77] ^ m[84] ^ m[85] ^ m[87] ^ m[90] ^ m[94] ^ m[99] ^ m[105] ^ m[112] ^ m[120] ^ m[121] ^ m[122] ^ m[123] ^ m[124] ^ m[126] ^ m[127] ^ m[128] ^ m[129] ^ m[131] ^ m[132] ^ m[133] ^ m[135] ^ m[136] ^ m[138] ^ m[141] ^ m[142] ^ m[143] ^ m[144] ^ m[146] ^ m[147] ^ m[148] ^ m[150] ^ m[151] ^ m[153] ^ m[156] ^ m[157] ^ m[158] ^ m[160] ^ m[161] ^ m[163] ^ m[166] ^ m[167] ^ m[169] ^ m[172] ^ m[176] ^ m[177] ^ m[178] ^ m[179] ^ m[181] ^ m[182] ^ m[183] ^ m[185] ^ m[186] ^ m[188] ^ m[191] ^ m[192] ^ m[193] ^ m[195] ^ m[196] ^ m[198] ^ m[201] ^ m[202] ^ m[204] ^ m[207] ^ m[211] ^ m[212] ^ m[213] ^ m[215] ^ m[216] ^ m[218] ^ m[221] ^ m[222] ^ m[224] ^ m[227] ^ m[231] ^ m[232] ^ m[234] ^ m[237] ^ m[241] ^ m[246] ^ m[247] ^ m[248] ^ m[249] ^ m[251] ^ m[252] ^ m[253] ^ m[255];
  end else if ((CodewordWidth == 523) && (MessageWidth == 512)) begin : gen_523_512
    `BR_ASSERT_STATIC(parity_width_matches_a, ParityWidth == 11)
    assign parity[0] = m[120] ^ m[121] ^ m[122] ^ m[123] ^ m[124] ^ m[125] ^ m[126] ^ m[127] ^ m[128] ^ m[129] ^ m[130] ^ m[131] ^ m[132] ^ m[133] ^ m[134] ^ m[135] ^ m[136] ^ m[137] ^ m[138] ^ m[139] ^ m[140] ^ m[141] ^ m[142] ^ m[143] ^ m[144] ^ m[145] ^ m[146] ^ m[147] ^ m[148] ^ m[149] ^ m[150] ^ m[151] ^ m[152] ^ m[153] ^ m[154] ^ m[155] ^ m[156] ^ m[157] ^ m[158] ^ m[159] ^ m[160] ^ m[161] ^ m[162] ^ m[163] ^ m[164] ^ m[417] ^ m[418] ^ m[419] ^ m[420] ^ m[421] ^ m[422] ^ m[423] ^ m[424] ^ m[425] ^ m[426] ^ m[427] ^ m[428] ^ m[429] ^ m[430] ^ m[431] ^ m[432] ^ m[433] ^ m[434] ^ m[435] ^ m[436] ^ m[437] ^ m[438] ^ m[439] ^ m[440] ^ m[441] ^ m[442] ^ m[443] ^ m[444] ^ m[445] ^ m[446] ^ m[447] ^ m[448] ^ m[449] ^ m[450] ^ m[451] ^ m[452] ^ m[453] ^ m[454] ^ m[455] ^ m[456] ^ m[457] ^ m[458] ^ m[459] ^ m[460] ^ m[461] ^ m[462] ^ m[463] ^ m[464] ^ m[465] ^ m[466] ^ m[467] ^ m[468] ^ m[469] ^ m[470] ^ m[471] ^ m[472] ^ m[473] ^ m[474] ^ m[475] ^ m[476] ^ m[477] ^ m[478] ^ m[479] ^ m[480] ^ m[481] ^ m[482] ^ m[483] ^ m[484] ^ m[485] ^ m[486] ^ m[487] ^ m[488] ^ m[489] ^ m[490] ^ m[491] ^ m[492] ^ m[493] ^ m[494] ^ m[495] ^ m[496] ^ m[497] ^ m[498] ^ m[499] ^ m[500] ^ m[501] ^ m[502] ^ m[503] ^ m[504] ^ m[505] ^ m[506] ^ m[507] ^ m[508] ^ m[509] ^ m[510] ^ m[511];
    assign parity[1] = m[84] ^ m[85] ^ m[86] ^ m[87] ^ m[88] ^ m[89] ^ m[90] ^ m[91] ^ m[92] ^ m[93] ^ m[94] ^ m[95] ^ m[96] ^ m[97] ^ m[98] ^ m[99] ^ m[100] ^ m[101] ^ m[102] ^ m[103] ^ m[104] ^ m[105] ^ m[106] ^ m[107] ^ m[108] ^ m[109] ^ m[110] ^ m[111] ^ m[112] ^ m[113] ^ m[114] ^ m[115] ^ m[116] ^ m[117] ^ m[118] ^ m[119] ^ m[156] ^ m[157] ^ m[158] ^ m[159] ^ m[160] ^ m[161] ^ m[162] ^ m[163] ^ m[164] ^ m[291] ^ m[292] ^ m[293] ^ m[294] ^ m[295] ^ m[296] ^ m[297] ^ m[298] ^ m[299] ^ m[300] ^ m[301] ^ m[302] ^ m[303] ^ m[304] ^ m[305] ^ m[306] ^ m[307] ^ m[308] ^ m[309] ^ m[310] ^ m[311] ^ m[312] ^ m[313] ^ m[314] ^ m[315] ^ m[316] ^ m[317] ^ m[318] ^ m[319] ^ m[320] ^ m[321] ^ m[322] ^ m[323] ^ m[324] ^ m[325] ^ m[326] ^ m[327] ^ m[328] ^ m[329] ^ m[330] ^ m[331] ^ m[332] ^ m[333] ^ m[334] ^ m[335] ^ m[336] ^ m[337] ^ m[338] ^ m[339] ^ m[340] ^ m[341] ^ m[342] ^ m[343] ^ m[344] ^ m[345] ^ m[346] ^ m[347] ^ m[348] ^ m[349] ^ m[350] ^ m[351] ^ m[352] ^ m[353] ^ m[354] ^ m[355] ^ m[356] ^ m[357] ^ m[358] ^ m[359] ^ m[360] ^ m[361] ^ m[362] ^ m[363] ^ m[364] ^ m[365] ^ m[366] ^ m[367] ^ m[368] ^ m[369] ^ m[370] ^ m[371] ^ m[372] ^ m[373] ^ m[374] ^ m[375] ^ m[376] ^ m[377] ^ m[378] ^ m[379] ^ m[380] ^ m[381] ^ m[382] ^ m[383] ^ m[384] ^ m[385] ^ m[386] ^ m[387] ^ m[388] ^ m[389] ^ m[390] ^ m[391] ^ m[392] ^ m[393] ^ m[394] ^ m[395] ^ m[396] ^ m[397] ^ m[398] ^ m[399] ^ m[400] ^ m[401] ^ m[402] ^ m[403] ^ m[404] ^ m[405] ^ m[406] ^ m[407] ^ m[408] ^ m[409] ^ m[410] ^ m[411] ^ m[412] ^ m[413] ^ m[414] ^ m[415] ^ m[416];
    assign parity[2] = m[56] ^ m[57] ^ m[58] ^ m[59] ^ m[60] ^ m[61] ^ m[62] ^ m[63] ^ m[64] ^ m[65] ^ m[66] ^ m[67] ^ m[68] ^ m[69] ^ m[70] ^ m[71] ^ m[72] ^ m[73] ^ m[74] ^ m[75] ^ m[76] ^ m[77] ^ m[78] ^ m[79] ^ m[80] ^ m[81] ^ m[82] ^ m[83] ^ m[112] ^ m[113] ^ m[114] ^ m[115] ^ m[116] ^ m[117] ^ m[118] ^ m[119] ^ m[148] ^ m[149] ^ m[150] ^ m[151] ^ m[152] ^ m[153] ^ m[154] ^ m[155] ^ m[164] ^ m[221] ^ m[222] ^ m[223] ^ m[224] ^ m[225] ^ m[226] ^ m[227] ^ m[228] ^ m[229] ^ m[230] ^ m[231] ^ m[232] ^ m[233] ^ m[234] ^ m[235] ^ m[236] ^ m[237] ^ m[238] ^ m[239] ^ m[240] ^ m[241] ^ m[242] ^ m[243] ^ m[244] ^ m[245] ^ m[246] ^ m[247] ^ m[248] ^ m[249] ^ m[250] ^ m[251] ^ m[252] ^ m[253] ^ m[254] ^ m[255] ^ m[256] ^ m[257] ^ m[258] ^ m[259] ^ m[260] ^ m[261] ^ m[262] ^ m[263] ^ m[264] ^ m[265] ^ m[266] ^ m[267] ^ m[268] ^ m[269] ^ m[270] ^ m[271] ^ m[272] ^ m[273] ^ m[274] ^ m[275] ^ m[276] ^ m[277] ^ m[278] ^ m[279] ^ m[280] ^ m[281] ^ m[282] ^ m[283] ^ m[284] ^ m[285] ^ m[286] ^ m[287] ^ m[288] ^ m[289] ^ m[290] ^ m[361] ^ m[362] ^ m[363] ^ m[364] ^ m[365] ^ m[366] ^ m[367] ^ m[368] ^ m[369] ^ m[370] ^ m[371] ^ m[372] ^ m[373] ^ m[374] ^ m[375] ^ m[376] ^ m[377] ^ m[378] ^ m[379] ^ m[380] ^ m[381] ^ m[382] ^ m[383] ^ m[384] ^ m[385] ^ m[386] ^ m[387] ^ m[388] ^ m[389] ^ m[390] ^ m[391] ^ m[392] ^ m[393] ^ m[394] ^ m[395] ^ m[396] ^ m[397] ^ m[398] ^ m[399] ^ m[400] ^ m[401] ^ m[402] ^ m[403] ^ m[404] ^ m[405] ^ m[406] ^ m[407] ^ m[408] ^ m[409] ^ m[410] ^ m[411] ^ m[412] ^ m[413] ^ m[414] ^ m[415] ^ m[416] ^ m[487] ^ m[488] ^ m[489] ^ m[490] ^ m[491] ^ m[492] ^ m[493] ^ m[494] ^ m[495] ^ m[496] ^ m[497] ^ m[498] ^ m[499] ^ m[500] ^ m[501] ^ m[502] ^ m[503] ^ m[504] ^ m[505] ^ m[506] ^ m[507] ^ m[508] ^ m[509] ^ m[510] ^ m[511];
    assign parity[3] = m[35] ^ m[36] ^ m[37] ^ m[38] ^ m[39] ^ m[40] ^ m[41] ^ m[42] ^ m[43] ^ m[44] ^ m[45] ^ m[46] ^ m[47] ^ m[48] ^ m[49] ^ m[50] ^ m[51] ^ m[52] ^ m[53] ^ m[54] ^ m[55] ^ m[77] ^ m[78] ^ m[79] ^ m[80] ^ m[81] ^ m[82] ^ m[83] ^ m[105] ^ m[106] ^ m[107] ^ m[108] ^ m[109] ^ m[110] ^ m[111] ^ m[119] ^ m[141] ^ m[142] ^ m[143] ^ m[144] ^ m[145] ^ m[146] ^ m[147] ^ m[155] ^ m[163] ^ m[186] ^ m[187] ^ m[188] ^ m[189] ^ m[190] ^ m[191] ^ m[192] ^ m[193] ^ m[194] ^ m[195] ^ m[196] ^ m[197] ^ m[198] ^ m[199] ^ m[200] ^ m[201] ^ m[202] ^ m[203] ^ m[204] ^ m[205] ^ m[206] ^ m[207] ^ m[208] ^ m[209] ^ m[210] ^ m[211] ^ m[212] ^ m[213] ^ m[214] ^ m[215] ^ m[216] ^ m[217] ^ m[218] ^ m[219] ^ m[220] ^ m[256] ^ m[257] ^ m[258] ^ m[259] ^ m[260] ^ m[261] ^ m[262] ^ m[263] ^ m[264] ^ m[265] ^ m[266] ^ m[267] ^ m[268] ^ m[269] ^ m[270] ^ m[271] ^ m[272] ^ m[273] ^ m[274] ^ m[275] ^ m[276] ^ m[277] ^ m[278] ^ m[279] ^ m[280] ^ m[281] ^ m[282] ^ m[283] ^ m[284] ^ m[285] ^ m[286] ^ m[287] ^ m[288] ^ m[289] ^ m[290] ^ m[326] ^ m[327] ^ m[328] ^ m[329] ^ m[330] ^ m[331] ^ m[332] ^ m[333] ^ m[334] ^ m[335] ^ m[336] ^ m[337] ^ m[338] ^ m[339] ^ m[340] ^ m[341] ^ m[342] ^ m[343] ^ m[344] ^ m[345] ^ m[346] ^ m[347] ^ m[348] ^ m[349] ^ m[350] ^ m[351] ^ m[352] ^ m[353] ^ m[354] ^ m[355] ^ m[356] ^ m[357] ^ m[358] ^ m[359] ^ m[360] ^ m[396] ^ m[397] ^ m[398] ^ m[399] ^ m[400] ^ m[401] ^ m[402] ^ m[403] ^ m[404] ^ m[405] ^ m[406] ^ m[407] ^ m[408] ^ m[409] ^ m[410] ^ m[411] ^ m[412] ^ m[413] ^ m[414] ^ m[415] ^ m[416] ^ m[452] ^ m[453] ^ m[454] ^ m[455] ^ m[456] ^ m[457] ^ m[458] ^ m[459] ^ m[460] ^ m[461] ^ m[462] ^ m[463] ^ m[464] ^ m[465] ^ m[466] ^ m[467] ^ m[468] ^ m[469] ^ m[470] ^ m[471] ^ m[472] ^ m[473] ^ m[474] ^ m[475] ^ m[476] ^ m[477] ^ m[478] ^ m[479] ^ m[480] ^ m[481] ^ m[482] ^ m[483] ^ m[484] ^ m[485] ^ m[486];
    assign parity[4] = m[20] ^ m[21] ^ m[22] ^ m[23] ^ m[24] ^ m[25] ^ m[26] ^ m[27] ^ m[28] ^ m[29] ^ m[30] ^ m[31] ^ m[32] ^ m[33] ^ m[34] ^ m[50] ^ m[51] ^ m[52] ^ m[53] ^ m[54] ^ m[55] ^ m[71] ^ m[72] ^ m[73] ^ m[74] ^ m[75] ^ m[76] ^ m[83] ^ m[99] ^ m[100] ^ m[101] ^ m[102] ^ m[103] ^ m[104] ^ m[111] ^ m[118] ^ m[135] ^ m[136] ^ m[137] ^ m[138] ^ m[139] ^ m[140] ^ m[147] ^ m[154] ^ m[162] ^ m[171] ^ m[172] ^ m[173] ^ m[174] ^ m[175] ^ m[176] ^ m[177] ^ m[178] ^ m[179] ^ m[180] ^ m[181] ^ m[182] ^ m[183] ^ m[184] ^ m[185] ^ m[201] ^ m[202] ^ m[203] ^ m[204] ^ m[205] ^ m[206] ^ m[207] ^ m[208] ^ m[209] ^ m[210] ^ m[211] ^ m[212] ^ m[213] ^ m[214] ^ m[215] ^ m[216] ^ m[217] ^ m[218] ^ m[219] ^ m[220] ^ m[236] ^ m[237] ^ m[238] ^ m[239] ^ m[240] ^ m[241] ^ m[242] ^ m[243] ^ m[244] ^ m[245] ^ m[246] ^ m[247] ^ m[248] ^ m[249] ^ m[250] ^ m[251] ^ m[252] ^ m[253] ^ m[254] ^ m[255] ^ m[276] ^ m[277] ^ m[278] ^ m[279] ^ m[280] ^ m[281] ^ m[282] ^ m[283] ^ m[284] ^ m[285] ^ m[286] ^ m[287] ^ m[288] ^ m[289] ^ m[290] ^ m[306] ^ m[307] ^ m[308] ^ m[309] ^ m[310] ^ m[311] ^ m[312] ^ m[313] ^ m[314] ^ m[315] ^ m[316] ^ m[317] ^ m[318] ^ m[319] ^ m[320] ^ m[321] ^ m[322] ^ m[323] ^ m[324] ^ m[325] ^ m[346] ^ m[347] ^ m[348] ^ m[349] ^ m[350] ^ m[351] ^ m[352] ^ m[353] ^ m[354] ^ m[355] ^ m[356] ^ m[357] ^ m[358] ^ m[359] ^ m[360] ^ m[381] ^ m[382] ^ m[383] ^ m[384] ^ m[385] ^ m[386] ^ m[387] ^ m[388] ^ m[389] ^ m[390] ^ m[391] ^ m[392] ^ m[393] ^ m[394] ^ m[395] ^ m[411] ^ m[412] ^ m[413] ^ m[414] ^ m[415] ^ m[416] ^ m[432] ^ m[433] ^ m[434] ^ m[435] ^ m[436] ^ m[437] ^ m[438] ^ m[439] ^ m[440] ^ m[441] ^ m[442] ^ m[443] ^ m[444] ^ m[445] ^ m[446] ^ m[447] ^ m[448] ^ m[449] ^ m[450] ^ m[451] ^ m[472] ^ m[473] ^ m[474] ^ m[475] ^ m[476] ^ m[477] ^ m[478] ^ m[479] ^ m[480] ^ m[481] ^ m[482] ^ m[483] ^ m[484] ^ m[485] ^ m[486] ^ m[507] ^ m[508] ^ m[509] ^ m[510] ^ m[511];
    assign parity[5] = m[10] ^ m[11] ^ m[12] ^ m[13] ^ m[14] ^ m[15] ^ m[16] ^ m[17] ^ m[18] ^ m[19] ^ m[30] ^ m[31] ^ m[32] ^ m[33] ^ m[34] ^ m[45] ^ m[46] ^ m[47] ^ m[48] ^ m[49] ^ m[55] ^ m[66] ^ m[67] ^ m[68] ^ m[69] ^ m[70] ^ m[76] ^ m[82] ^ m[94] ^ m[95] ^ m[96] ^ m[97] ^ m[98] ^ m[104] ^ m[110] ^ m[117] ^ m[130] ^ m[131] ^ m[132] ^ m[133] ^ m[134] ^ m[140] ^ m[146] ^ m[153] ^ m[161] ^ m[166] ^ m[167] ^ m[168] ^ m[169] ^ m[170] ^ m[176] ^ m[177] ^ m[178] ^ m[179] ^ m[180] ^ m[181] ^ m[182] ^ m[183] ^ m[184] ^ m[185] ^ m[191] ^ m[192] ^ m[193] ^ m[194] ^ m[195] ^ m[196] ^ m[197] ^ m[198] ^ m[199] ^ m[200] ^ m[211] ^ m[212] ^ m[213] ^ m[214] ^ m[215] ^ m[216] ^ m[217] ^ m[218] ^ m[219] ^ m[220] ^ m[226] ^ m[227] ^ m[228] ^ m[229] ^ m[230] ^ m[231] ^ m[232] ^ m[233] ^ m[234] ^ m[235] ^ m[246] ^ m[247] ^ m[248] ^ m[249] ^ m[250] ^ m[251] ^ m[252] ^ m[253] ^ m[254] ^ m[255] ^ m[266] ^ m[267] ^ m[268] ^ m[269] ^ m[270] ^ m[271] ^ m[272] ^ m[273] ^ m[274] ^ m[275] ^ m[286] ^ m[287] ^ m[288] ^ m[289] ^ m[290] ^ m[296] ^ m[297] ^ m[298] ^ m[299] ^ m[300] ^ m[301] ^ m[302] ^ m[303] ^ m[304] ^ m[305] ^ m[316] ^ m[317] ^ m[318] ^ m[319] ^ m[320] ^ m[321] ^ m[322] ^ m[323] ^ m[324] ^ m[325] ^ m[336] ^ m[337] ^ m[338] ^ m[339] ^ m[340] ^ m[341] ^ m[342] ^ m[343] ^ m[344] ^ m[345] ^ m[356] ^ m[357] ^ m[358] ^ m[359] ^ m[360] ^ m[371] ^ m[372] ^ m[373] ^ m[374] ^ m[375] ^ m[376] ^ m[377] ^ m[378] ^ m[379] ^ m[380] ^ m[391] ^ m[392] ^ m[393] ^ m[394] ^ m[395] ^ m[406] ^ m[407] ^ m[408] ^ m[409] ^ m[410] ^ m[416] ^ m[422] ^ m[423] ^ m[424] ^ m[425] ^ m[426] ^ m[427] ^ m[428] ^ m[429] ^ m[430] ^ m[431] ^ m[442] ^ m[443] ^ m[444] ^ m[445] ^ m[446] ^ m[447] ^ m[448] ^ m[449] ^ m[450] ^ m[451] ^ m[462] ^ m[463] ^ m[464] ^ m[465] ^ m[466] ^ m[467] ^ m[468] ^ m[469] ^ m[470] ^ m[471] ^ m[482] ^ m[483] ^ m[484] ^ m[485] ^ m[486] ^ m[497] ^ m[498] ^ m[499] ^ m[500] ^ m[501] ^ m[502] ^ m[503] ^ m[504] ^ m[505] ^ m[506];
    assign parity[6] = m[4] ^ m[5] ^ m[6] ^ m[7] ^ m[8] ^ m[9] ^ m[16] ^ m[17] ^ m[18] ^ m[19] ^ m[26] ^ m[27] ^ m[28] ^ m[29] ^ m[34] ^ m[41] ^ m[42] ^ m[43] ^ m[44] ^ m[49] ^ m[54] ^ m[62] ^ m[63] ^ m[64] ^ m[65] ^ m[70] ^ m[75] ^ m[81] ^ m[90] ^ m[91] ^ m[92] ^ m[93] ^ m[98] ^ m[103] ^ m[109] ^ m[116] ^ m[126] ^ m[127] ^ m[128] ^ m[129] ^ m[134] ^ m[139] ^ m[145] ^ m[152] ^ m[160] ^ m[165] ^ m[167] ^ m[168] ^ m[169] ^ m[170] ^ m[172] ^ m[173] ^ m[174] ^ m[175] ^ m[180] ^ m[181] ^ m[182] ^ m[183] ^ m[184] ^ m[185] ^ m[187] ^ m[188] ^ m[189] ^ m[190] ^ m[195] ^ m[196] ^ m[197] ^ m[198] ^ m[199] ^ m[200] ^ m[205] ^ m[206] ^ m[207] ^ m[208] ^ m[209] ^ m[210] ^ m[217] ^ m[218] ^ m[219] ^ m[220] ^ m[222] ^ m[223] ^ m[224] ^ m[225] ^ m[230] ^ m[231] ^ m[232] ^ m[233] ^ m[234] ^ m[235] ^ m[240] ^ m[241] ^ m[242] ^ m[243] ^ m[244] ^ m[245] ^ m[252] ^ m[253] ^ m[254] ^ m[255] ^ m[260] ^ m[261] ^ m[262] ^ m[263] ^ m[264] ^ m[265] ^ m[272] ^ m[273] ^ m[274] ^ m[275] ^ m[282] ^ m[283] ^ m[284] ^ m[285] ^ m[290] ^ m[292] ^ m[293] ^ m[294] ^ m[295] ^ m[300] ^ m[301] ^ m[302] ^ m[303] ^ m[304] ^ m[305] ^ m[310] ^ m[311] ^ m[312] ^ m[313] ^ m[314] ^ m[315] ^ m[322] ^ m[323] ^ m[324] ^ m[325] ^ m[330] ^ m[331] ^ m[332] ^ m[333] ^ m[334] ^ m[335] ^ m[342] ^ m[343] ^ m[344] ^ m[345] ^ m[352] ^ m[353] ^ m[354] ^ m[355] ^ m[360] ^ m[365] ^ m[366] ^ m[367] ^ m[368] ^ m[369] ^ m[370] ^ m[377] ^ m[378] ^ m[379] ^ m[380] ^ m[387] ^ m[388] ^ m[389] ^ m[390] ^ m[395] ^ m[402] ^ m[403] ^ m[404] ^ m[405] ^ m[410] ^ m[415] ^ m[418] ^ m[419] ^ m[420] ^ m[421] ^ m[426] ^ m[427] ^ m[428] ^ m[429] ^ m[430] ^ m[431] ^ m[436] ^ m[437] ^ m[438] ^ m[439] ^ m[440] ^ m[441] ^ m[448] ^ m[449] ^ m[450] ^ m[451] ^ m[456] ^ m[457] ^ m[458] ^ m[459] ^ m[460] ^ m[461] ^ m[468] ^ m[469] ^ m[470] ^ m[471] ^ m[478] ^ m[479] ^ m[480] ^ m[481] ^ m[486] ^ m[491] ^ m[492] ^ m[493] ^ m[494] ^ m[495] ^ m[496] ^ m[503] ^ m[504] ^ m[505] ^ m[506];
    assign parity[7] = m[1] ^ m[2] ^ m[3] ^ m[7] ^ m[8] ^ m[9] ^ m[13] ^ m[14] ^ m[15] ^ m[19] ^ m[23] ^ m[24] ^ m[25] ^ m[29] ^ m[33] ^ m[38] ^ m[39] ^ m[40] ^ m[44] ^ m[48] ^ m[53] ^ m[59] ^ m[60] ^ m[61] ^ m[65] ^ m[69] ^ m[74] ^ m[80] ^ m[87] ^ m[88] ^ m[89] ^ m[93] ^ m[97] ^ m[102] ^ m[108] ^ m[115] ^ m[123] ^ m[124] ^ m[125] ^ m[129] ^ m[133] ^ m[138] ^ m[144] ^ m[151] ^ m[159] ^ m[165] ^ m[166] ^ m[168] ^ m[169] ^ m[170] ^ m[171] ^ m[173] ^ m[174] ^ m[175] ^ m[177] ^ m[178] ^ m[179] ^ m[183] ^ m[184] ^ m[185] ^ m[186] ^ m[188] ^ m[189] ^ m[190] ^ m[192] ^ m[193] ^ m[194] ^ m[198] ^ m[199] ^ m[200] ^ m[202] ^ m[203] ^ m[204] ^ m[208] ^ m[209] ^ m[210] ^ m[214] ^ m[215] ^ m[216] ^ m[220] ^ m[221] ^ m[223] ^ m[224] ^ m[225] ^ m[227] ^ m[228] ^ m[229] ^ m[233] ^ m[234] ^ m[235] ^ m[237] ^ m[238] ^ m[239] ^ m[243] ^ m[244] ^ m[245] ^ m[249] ^ m[250] ^ m[251] ^ m[255] ^ m[257] ^ m[258] ^ m[259] ^ m[263] ^ m[264] ^ m[265] ^ m[269] ^ m[270] ^ m[271] ^ m[275] ^ m[279] ^ m[280] ^ m[281] ^ m[285] ^ m[289] ^ m[291] ^ m[293] ^ m[294] ^ m[295] ^ m[297] ^ m[298] ^ m[299] ^ m[303] ^ m[304] ^ m[305] ^ m[307] ^ m[308] ^ m[309] ^ m[313] ^ m[314] ^ m[315] ^ m[319] ^ m[320] ^ m[321] ^ m[325] ^ m[327] ^ m[328] ^ m[329] ^ m[333] ^ m[334] ^ m[335] ^ m[339] ^ m[340] ^ m[341] ^ m[345] ^ m[349] ^ m[350] ^ m[351] ^ m[355] ^ m[359] ^ m[362] ^ m[363] ^ m[364] ^ m[368] ^ m[369] ^ m[370] ^ m[374] ^ m[375] ^ m[376] ^ m[380] ^ m[384] ^ m[385] ^ m[386] ^ m[390] ^ m[394] ^ m[399] ^ m[400] ^ m[401] ^ m[405] ^ m[409] ^ m[414] ^ m[417] ^ m[419] ^ m[420] ^ m[421] ^ m[423] ^ m[424] ^ m[425] ^ m[429] ^ m[430] ^ m[431] ^ m[433] ^ m[434] ^ m[435] ^ m[439] ^ m[440] ^ m[441] ^ m[445] ^ m[446] ^ m[447] ^ m[451] ^ m[453] ^ m[454] ^ m[455] ^ m[459] ^ m[460] ^ m[461] ^ m[465] ^ m[466] ^ m[467] ^ m[471] ^ m[475] ^ m[476] ^ m[477] ^ m[481] ^ m[485] ^ m[488] ^ m[489] ^ m[490] ^ m[494] ^ m[495] ^ m[496] ^ m[500] ^ m[501] ^ m[502] ^ m[506] ^ m[510] ^ m[511];
    assign parity[8] = m[0] ^ m[2] ^ m[3] ^ m[5] ^ m[6] ^ m[9] ^ m[11] ^ m[12] ^ m[15] ^ m[18] ^ m[21] ^ m[22] ^ m[25] ^ m[28] ^ m[32] ^ m[36] ^ m[37] ^ m[40] ^ m[43] ^ m[47] ^ m[52] ^ m[57] ^ m[58] ^ m[61] ^ m[64] ^ m[68] ^ m[73] ^ m[79] ^ m[85] ^ m[86] ^ m[89] ^ m[92] ^ m[96] ^ m[101] ^ m[107] ^ m[114] ^ m[121] ^ m[122] ^ m[125] ^ m[128] ^ m[132] ^ m[137] ^ m[143] ^ m[150] ^ m[158] ^ m[165] ^ m[166] ^ m[167] ^ m[169] ^ m[170] ^ m[171] ^ m[172] ^ m[174] ^ m[175] ^ m[176] ^ m[178] ^ m[179] ^ m[181] ^ m[182] ^ m[185] ^ m[186] ^ m[187] ^ m[189] ^ m[190] ^ m[191] ^ m[193] ^ m[194] ^ m[196] ^ m[197] ^ m[200] ^ m[201] ^ m[203] ^ m[204] ^ m[206] ^ m[207] ^ m[210] ^ m[212] ^ m[213] ^ m[216] ^ m[219] ^ m[221] ^ m[222] ^ m[224] ^ m[225] ^ m[226] ^ m[228] ^ m[229] ^ m[231] ^ m[232] ^ m[235] ^ m[236] ^ m[238] ^ m[239] ^ m[241] ^ m[242] ^ m[245] ^ m[247] ^ m[248] ^ m[251] ^ m[254] ^ m[256] ^ m[258] ^ m[259] ^ m[261] ^ m[262] ^ m[265] ^ m[267] ^ m[268] ^ m[271] ^ m[274] ^ m[277] ^ m[278] ^ m[281] ^ m[284] ^ m[288] ^ m[291] ^ m[292] ^ m[294] ^ m[295] ^ m[296] ^ m[298] ^ m[299] ^ m[301] ^ m[302] ^ m[305] ^ m[306] ^ m[308] ^ m[309] ^ m[311] ^ m[312] ^ m[315] ^ m[317] ^ m[318] ^ m[321] ^ m[324] ^ m[326] ^ m[328] ^ m[329] ^ m[331] ^ m[332] ^ m[335] ^ m[337] ^ m[338] ^ m[341] ^ m[344] ^ m[347] ^ m[348] ^ m[351] ^ m[354] ^ m[358] ^ m[361] ^ m[363] ^ m[364] ^ m[366] ^ m[367] ^ m[370] ^ m[372] ^ m[373] ^ m[376] ^ m[379] ^ m[382] ^ m[383] ^ m[386] ^ m[389] ^ m[393] ^ m[397] ^ m[398] ^ m[401] ^ m[404] ^ m[408] ^ m[413] ^ m[417] ^ m[418] ^ m[420] ^ m[421] ^ m[422] ^ m[424] ^ m[425] ^ m[427] ^ m[428] ^ m[431] ^ m[432] ^ m[434] ^ m[435] ^ m[437] ^ m[438] ^ m[441] ^ m[443] ^ m[444] ^ m[447] ^ m[450] ^ m[452] ^ m[454] ^ m[455] ^ m[457] ^ m[458] ^ m[461] ^ m[463] ^ m[464] ^ m[467] ^ m[470] ^ m[473] ^ m[474] ^ m[477] ^ m[480] ^ m[484] ^ m[487] ^ m[489] ^ m[490] ^ m[492] ^ m[493] ^ m[496] ^ m[498] ^ m[499] ^ m[502] ^ m[505] ^ m[508] ^ m[509];
    assign parity[9] = m[0] ^ m[1] ^ m[3] ^ m[4] ^ m[6] ^ m[8] ^ m[10] ^ m[12] ^ m[14] ^ m[17] ^ m[20] ^ m[22] ^ m[24] ^ m[27] ^ m[31] ^ m[35] ^ m[37] ^ m[39] ^ m[42] ^ m[46] ^ m[51] ^ m[56] ^ m[58] ^ m[60] ^ m[63] ^ m[67] ^ m[72] ^ m[78] ^ m[84] ^ m[86] ^ m[88] ^ m[91] ^ m[95] ^ m[100] ^ m[106] ^ m[113] ^ m[120] ^ m[122] ^ m[124] ^ m[127] ^ m[131] ^ m[136] ^ m[142] ^ m[149] ^ m[157] ^ m[165] ^ m[166] ^ m[167] ^ m[168] ^ m[170] ^ m[171] ^ m[172] ^ m[173] ^ m[175] ^ m[176] ^ m[177] ^ m[179] ^ m[180] ^ m[182] ^ m[184] ^ m[186] ^ m[187] ^ m[188] ^ m[190] ^ m[191] ^ m[192] ^ m[194] ^ m[195] ^ m[197] ^ m[199] ^ m[201] ^ m[202] ^ m[204] ^ m[205] ^ m[207] ^ m[209] ^ m[211] ^ m[213] ^ m[215] ^ m[218] ^ m[221] ^ m[222] ^ m[223] ^ m[225] ^ m[226] ^ m[227] ^ m[229] ^ m[230] ^ m[232] ^ m[234] ^ m[236] ^ m[237] ^ m[239] ^ m[240] ^ m[242] ^ m[244] ^ m[246] ^ m[248] ^ m[250] ^ m[253] ^ m[256] ^ m[257] ^ m[259] ^ m[260] ^ m[262] ^ m[264] ^ m[266] ^ m[268] ^ m[270] ^ m[273] ^ m[276] ^ m[278] ^ m[280] ^ m[283] ^ m[287] ^ m[291] ^ m[292] ^ m[293] ^ m[295] ^ m[296] ^ m[297] ^ m[299] ^ m[300] ^ m[302] ^ m[304] ^ m[306] ^ m[307] ^ m[309] ^ m[310] ^ m[312] ^ m[314] ^ m[316] ^ m[318] ^ m[320] ^ m[323] ^ m[326] ^ m[327] ^ m[329] ^ m[330] ^ m[332] ^ m[334] ^ m[336] ^ m[338] ^ m[340] ^ m[343] ^ m[346] ^ m[348] ^ m[350] ^ m[353] ^ m[357] ^ m[361] ^ m[362] ^ m[364] ^ m[365] ^ m[367] ^ m[369] ^ m[371] ^ m[373] ^ m[375] ^ m[378] ^ m[381] ^ m[383] ^ m[385] ^ m[388] ^ m[392] ^ m[396] ^ m[398] ^ m[400] ^ m[403] ^ m[407] ^ m[412] ^ m[417] ^ m[418] ^ m[419] ^ m[421] ^ m[422] ^ m[423] ^ m[425] ^ m[426] ^ m[428] ^ m[430] ^ m[432] ^ m[433] ^ m[435] ^ m[436] ^ m[438] ^ m[440] ^ m[442] ^ m[444] ^ m[446] ^ m[449] ^ m[452] ^ m[453] ^ m[455] ^ m[456] ^ m[458] ^ m[460] ^ m[462] ^ m[464] ^ m[466] ^ m[469] ^ m[472] ^ m[474] ^ m[476] ^ m[479] ^ m[483] ^ m[487] ^ m[488] ^ m[490] ^ m[491] ^ m[493] ^ m[495] ^ m[497] ^ m[499] ^ m[501] ^ m[504] ^ m[507] ^ m[509] ^ m[511];
    assign parity[10] = m[0] ^ m[1] ^ m[2] ^ m[4] ^ m[5] ^ m[7] ^ m[10] ^ m[11] ^ m[13] ^ m[16] ^ m[20] ^ m[21] ^ m[23] ^ m[26] ^ m[30] ^ m[35] ^ m[36] ^ m[38] ^ m[41] ^ m[45] ^ m[50] ^ m[56] ^ m[57] ^ m[59] ^ m[62] ^ m[66] ^ m[71] ^ m[77] ^ m[84] ^ m[85] ^ m[87] ^ m[90] ^ m[94] ^ m[99] ^ m[105] ^ m[112] ^ m[120] ^ m[121] ^ m[123] ^ m[126] ^ m[130] ^ m[135] ^ m[141] ^ m[148] ^ m[156] ^ m[165] ^ m[166] ^ m[167] ^ m[168] ^ m[169] ^ m[171] ^ m[172] ^ m[173] ^ m[174] ^ m[176] ^ m[177] ^ m[178] ^ m[180] ^ m[181] ^ m[183] ^ m[186] ^ m[187] ^ m[188] ^ m[189] ^ m[191] ^ m[192] ^ m[193] ^ m[195] ^ m[196] ^ m[198] ^ m[201] ^ m[202] ^ m[203] ^ m[205] ^ m[206] ^ m[208] ^ m[211] ^ m[212] ^ m[214] ^ m[217] ^ m[221] ^ m[222] ^ m[223] ^ m[224] ^ m[226] ^ m[227] ^ m[228] ^ m[230] ^ m[231] ^ m[233] ^ m[236] ^ m[237] ^ m[238] ^ m[240] ^ m[241] ^ m[243] ^ m[246] ^ m[247] ^ m[249] ^ m[252] ^ m[256] ^ m[257] ^ m[258] ^ m[260] ^ m[261] ^ m[263] ^ m[266] ^ m[267] ^ m[269] ^ m[272] ^ m[276] ^ m[277] ^ m[279] ^ m[282] ^ m[286] ^ m[291] ^ m[292] ^ m[293] ^ m[294] ^ m[296] ^ m[297] ^ m[298] ^ m[300] ^ m[301] ^ m[303] ^ m[306] ^ m[307] ^ m[308] ^ m[310] ^ m[311] ^ m[313] ^ m[316] ^ m[317] ^ m[319] ^ m[322] ^ m[326] ^ m[327] ^ m[328] ^ m[330] ^ m[331] ^ m[333] ^ m[336] ^ m[337] ^ m[339] ^ m[342] ^ m[346] ^ m[347] ^ m[349] ^ m[352] ^ m[356] ^ m[361] ^ m[362] ^ m[363] ^ m[365] ^ m[366] ^ m[368] ^ m[371] ^ m[372] ^ m[374] ^ m[377] ^ m[381] ^ m[382] ^ m[384] ^ m[387] ^ m[391] ^ m[396] ^ m[397] ^ m[399] ^ m[402] ^ m[406] ^ m[411] ^ m[417] ^ m[418] ^ m[419] ^ m[420] ^ m[422] ^ m[423] ^ m[424] ^ m[426] ^ m[427] ^ m[429] ^ m[432] ^ m[433] ^ m[434] ^ m[436] ^ m[437] ^ m[439] ^ m[442] ^ m[443] ^ m[445] ^ m[448] ^ m[452] ^ m[453] ^ m[454] ^ m[456] ^ m[457] ^ m[459] ^ m[462] ^ m[463] ^ m[465] ^ m[468] ^ m[472] ^ m[473] ^ m[475] ^ m[478] ^ m[482] ^ m[487] ^ m[488] ^ m[489] ^ m[491] ^ m[492] ^ m[494] ^ m[497] ^ m[498] ^ m[500] ^ m[503] ^ m[507] ^ m[508] ^ m[510];
  end else if ((CodewordWidth == 1036) && (MessageWidth == 1024)) begin : gen_1036_1024
    `BR_ASSERT_STATIC(parity_width_matches_a, ParityWidth == 12)
    assign parity[0] = m[165] ^ m[166] ^ m[167] ^ m[168] ^ m[169] ^ m[170] ^ m[171] ^ m[172] ^ m[173] ^ m[174] ^ m[175] ^ m[176] ^ m[177] ^ m[178] ^ m[179] ^ m[180] ^ m[181] ^ m[182] ^ m[183] ^ m[184] ^ m[185] ^ m[186] ^ m[187] ^ m[188] ^ m[189] ^ m[190] ^ m[191] ^ m[192] ^ m[193] ^ m[194] ^ m[195] ^ m[196] ^ m[197] ^ m[198] ^ m[199] ^ m[200] ^ m[201] ^ m[202] ^ m[203] ^ m[204] ^ m[205] ^ m[206] ^ m[207] ^ m[208] ^ m[209] ^ m[210] ^ m[211] ^ m[212] ^ m[213] ^ m[214] ^ m[215] ^ m[216] ^ m[217] ^ m[218] ^ m[219] ^ m[682] ^ m[683] ^ m[684] ^ m[685] ^ m[686] ^ m[687] ^ m[688] ^ m[689] ^ m[690] ^ m[691] ^ m[692] ^ m[693] ^ m[694] ^ m[695] ^ m[696] ^ m[697] ^ m[698] ^ m[699] ^ m[700] ^ m[701] ^ m[702] ^ m[703] ^ m[704] ^ m[705] ^ m[706] ^ m[707] ^ m[708] ^ m[709] ^ m[710] ^ m[711] ^ m[712] ^ m[713] ^ m[714] ^ m[715] ^ m[716] ^ m[717] ^ m[718] ^ m[719] ^ m[720] ^ m[721] ^ m[722] ^ m[723] ^ m[724] ^ m[725] ^ m[726] ^ m[727] ^ m[728] ^ m[729] ^ m[730] ^ m[731] ^ m[732] ^ m[733] ^ m[734] ^ m[735] ^ m[736] ^ m[737] ^ m[738] ^ m[739] ^ m[740] ^ m[741] ^ m[742] ^ m[743] ^ m[744] ^ m[745] ^ m[746] ^ m[747] ^ m[748] ^ m[749] ^ m[750] ^ m[751] ^ m[752] ^ m[753] ^ m[754] ^ m[755] ^ m[756] ^ m[757] ^ m[758] ^ m[759] ^ m[760] ^ m[761] ^ m[762] ^ m[763] ^ m[764] ^ m[765] ^ m[766] ^ m[767] ^ m[768] ^ m[769] ^ m[770] ^ m[771] ^ m[772] ^ m[773] ^ m[774] ^ m[775] ^ m[776] ^ m[777] ^ m[778] ^ m[779] ^ m[780] ^ m[781] ^ m[782] ^ m[783] ^ m[784] ^ m[785] ^ m[786] ^ m[787] ^ m[788] ^ m[789] ^ m[790] ^ m[791] ^ m[792] ^ m[793] ^ m[794] ^ m[795] ^ m[796] ^ m[797] ^ m[798] ^ m[799] ^ m[800] ^ m[801] ^ m[802] ^ m[803] ^ m[804] ^ m[805] ^ m[806] ^ m[807] ^ m[808] ^ m[809] ^ m[810] ^ m[811] ^ m[812] ^ m[813] ^ m[814] ^ m[815] ^ m[816] ^ m[817] ^ m[818] ^ m[819] ^ m[820] ^ m[821] ^ m[822] ^ m[823] ^ m[824] ^ m[825] ^ m[826] ^ m[827] ^ m[828] ^ m[829] ^ m[830] ^ m[831] ^ m[832] ^ m[833] ^ m[834] ^ m[835] ^ m[836] ^ m[837] ^ m[838] ^ m[839] ^ m[840] ^ m[841] ^ m[842] ^ m[843] ^ m[844] ^ m[845] ^ m[846] ^ m[847] ^ m[848] ^ m[849] ^ m[850] ^ m[851] ^ m[852] ^ m[853] ^ m[854] ^ m[855] ^ m[856] ^ m[857] ^ m[858] ^ m[859] ^ m[860] ^ m[861] ^ m[862] ^ m[863] ^ m[864] ^ m[865] ^ m[866] ^ m[867] ^ m[868] ^ m[869] ^ m[870] ^ m[871] ^ m[872] ^ m[873] ^ m[874] ^ m[875] ^ m[876] ^ m[877] ^ m[878] ^ m[879] ^ m[880] ^ m[881] ^ m[882] ^ m[883] ^ m[884] ^ m[885] ^ m[886] ^ m[887] ^ m[888] ^ m[889] ^ m[890] ^ m[891] ^ m[892] ^ m[893] ^ m[894] ^ m[895] ^ m[896] ^ m[897] ^ m[898] ^ m[899] ^ m[900] ^ m[901] ^ m[902] ^ m[903] ^ m[904] ^ m[905] ^ m[906] ^ m[907] ^ m[908] ^ m[909] ^ m[910] ^ m[911] ^ m[912] ^ m[913] ^ m[914] ^ m[915] ^ m[916] ^ m[917] ^ m[918] ^ m[919] ^ m[920] ^ m[921] ^ m[922] ^ m[923] ^ m[924] ^ m[925] ^ m[926] ^ m[927] ^ m[928] ^ m[929] ^ m[930] ^ m[931] ^ m[932] ^ m[933] ^ m[934] ^ m[935] ^ m[936] ^ m[937] ^ m[938] ^ m[939] ^ m[940] ^ m[941] ^ m[942] ^ m[943] ^ m[944] ^ m[945] ^ m[946] ^ m[947] ^ m[948] ^ m[949] ^ m[950] ^ m[951] ^ m[952] ^ m[953] ^ m[954] ^ m[955] ^ m[956] ^ m[957] ^ m[958] ^ m[959] ^ m[960] ^ m[961] ^ m[962] ^ m[963] ^ m[964] ^ m[965] ^ m[966] ^ m[967] ^ m[968] ^ m[969] ^ m[970] ^ m[971] ^ m[972] ^ m[973] ^ m[974] ^ m[975] ^ m[976] ^ m[977] ^ m[978] ^ m[979] ^ m[980] ^ m[981] ^ m[982] ^ m[983] ^ m[984] ^ m[985] ^ m[986] ^ m[987] ^ m[988] ^ m[989] ^ m[990] ^ m[991] ^ m[992] ^ m[993] ^ m[994] ^ m[995] ^ m[996] ^ m[997] ^ m[998] ^ m[999] ^ m[1000] ^ m[1001] ^ m[1002] ^ m[1003] ^ m[1004] ^ m[1005] ^ m[1006] ^ m[1007] ^ m[1008] ^ m[1009] ^ m[1010] ^ m[1011];
    assign parity[1] = m[120] ^ m[121] ^ m[122] ^ m[123] ^ m[124] ^ m[125] ^ m[126] ^ m[127] ^ m[128] ^ m[129] ^ m[130] ^ m[131] ^ m[132] ^ m[133] ^ m[134] ^ m[135] ^ m[136] ^ m[137] ^ m[138] ^ m[139] ^ m[140] ^ m[141] ^ m[142] ^ m[143] ^ m[144] ^ m[145] ^ m[146] ^ m[147] ^ m[148] ^ m[149] ^ m[150] ^ m[151] ^ m[152] ^ m[153] ^ m[154] ^ m[155] ^ m[156] ^ m[157] ^ m[158] ^ m[159] ^ m[160] ^ m[161] ^ m[162] ^ m[163] ^ m[164] ^ m[210] ^ m[211] ^ m[212] ^ m[213] ^ m[214] ^ m[215] ^ m[216] ^ m[217] ^ m[218] ^ m[219] ^ m[472] ^ m[473] ^ m[474] ^ m[475] ^ m[476] ^ m[477] ^ m[478] ^ m[479] ^ m[480] ^ m[481] ^ m[482] ^ m[483] ^ m[484] ^ m[485] ^ m[486] ^ m[487] ^ m[488] ^ m[489] ^ m[490] ^ m[491] ^ m[492] ^ m[493] ^ m[494] ^ m[495] ^ m[496] ^ m[497] ^ m[498] ^ m[499] ^ m[500] ^ m[501] ^ m[502] ^ m[503] ^ m[504] ^ m[505] ^ m[506] ^ m[507] ^ m[508] ^ m[509] ^ m[510] ^ m[511] ^ m[512] ^ m[513] ^ m[514] ^ m[515] ^ m[516] ^ m[517] ^ m[518] ^ m[519] ^ m[520] ^ m[521] ^ m[522] ^ m[523] ^ m[524] ^ m[525] ^ m[526] ^ m[527] ^ m[528] ^ m[529] ^ m[530] ^ m[531] ^ m[532] ^ m[533] ^ m[534] ^ m[535] ^ m[536] ^ m[537] ^ m[538] ^ m[539] ^ m[540] ^ m[541] ^ m[542] ^ m[543] ^ m[544] ^ m[545] ^ m[546] ^ m[547] ^ m[548] ^ m[549] ^ m[550] ^ m[551] ^ m[552] ^ m[553] ^ m[554] ^ m[555] ^ m[556] ^ m[557] ^ m[558] ^ m[559] ^ m[560] ^ m[561] ^ m[562] ^ m[563] ^ m[564] ^ m[565] ^ m[566] ^ m[567] ^ m[568] ^ m[569] ^ m[570] ^ m[571] ^ m[572] ^ m[573] ^ m[574] ^ m[575] ^ m[576] ^ m[577] ^ m[578] ^ m[579] ^ m[580] ^ m[581] ^ m[582] ^ m[583] ^ m[584] ^ m[585] ^ m[586] ^ m[587] ^ m[588] ^ m[589] ^ m[590] ^ m[591] ^ m[592] ^ m[593] ^ m[594] ^ m[595] ^ m[596] ^ m[597] ^ m[598] ^ m[599] ^ m[600] ^ m[601] ^ m[602] ^ m[603] ^ m[604] ^ m[605] ^ m[606] ^ m[607] ^ m[608] ^ m[609] ^ m[610] ^ m[611] ^ m[612] ^ m[613] ^ m[614] ^ m[615] ^ m[616] ^ m[617] ^ m[618] ^ m[619] ^ m[620] ^ m[621] ^ m[622] ^ m[623] ^ m[624] ^ m[625] ^ m[626] ^ m[627] ^ m[628] ^ m[629] ^ m[630] ^ m[631] ^ m[632] ^ m[633] ^ m[634] ^ m[635] ^ m[636] ^ m[637] ^ m[638] ^ m[639] ^ m[640] ^ m[641] ^ m[642] ^ m[643] ^ m[644] ^ m[645] ^ m[646] ^ m[647] ^ m[648] ^ m[649] ^ m[650] ^ m[651] ^ m[652] ^ m[653] ^ m[654] ^ m[655] ^ m[656] ^ m[657] ^ m[658] ^ m[659] ^ m[660] ^ m[661] ^ m[662] ^ m[663] ^ m[664] ^ m[665] ^ m[666] ^ m[667] ^ m[668] ^ m[669] ^ m[670] ^ m[671] ^ m[672] ^ m[673] ^ m[674] ^ m[675] ^ m[676] ^ m[677] ^ m[678] ^ m[679] ^ m[680] ^ m[681] ^ m[892] ^ m[893] ^ m[894] ^ m[895] ^ m[896] ^ m[897] ^ m[898] ^ m[899] ^ m[900] ^ m[901] ^ m[902] ^ m[903] ^ m[904] ^ m[905] ^ m[906] ^ m[907] ^ m[908] ^ m[909] ^ m[910] ^ m[911] ^ m[912] ^ m[913] ^ m[914] ^ m[915] ^ m[916] ^ m[917] ^ m[918] ^ m[919] ^ m[920] ^ m[921] ^ m[922] ^ m[923] ^ m[924] ^ m[925] ^ m[926] ^ m[927] ^ m[928] ^ m[929] ^ m[930] ^ m[931] ^ m[932] ^ m[933] ^ m[934] ^ m[935] ^ m[936] ^ m[937] ^ m[938] ^ m[939] ^ m[940] ^ m[941] ^ m[942] ^ m[943] ^ m[944] ^ m[945] ^ m[946] ^ m[947] ^ m[948] ^ m[949] ^ m[950] ^ m[951] ^ m[952] ^ m[953] ^ m[954] ^ m[955] ^ m[956] ^ m[957] ^ m[958] ^ m[959] ^ m[960] ^ m[961] ^ m[962] ^ m[963] ^ m[964] ^ m[965] ^ m[966] ^ m[967] ^ m[968] ^ m[969] ^ m[970] ^ m[971] ^ m[972] ^ m[973] ^ m[974] ^ m[975] ^ m[976] ^ m[977] ^ m[978] ^ m[979] ^ m[980] ^ m[981] ^ m[982] ^ m[983] ^ m[984] ^ m[985] ^ m[986] ^ m[987] ^ m[988] ^ m[989] ^ m[990] ^ m[991] ^ m[992] ^ m[993] ^ m[994] ^ m[995] ^ m[996] ^ m[997] ^ m[998] ^ m[999] ^ m[1000] ^ m[1001] ^ m[1002] ^ m[1003] ^ m[1004] ^ m[1005] ^ m[1006] ^ m[1007] ^ m[1008] ^ m[1009] ^ m[1010] ^ m[1011];
    assign parity[2] = m[84] ^ m[85] ^ m[86] ^ m[87] ^ m[88] ^ m[89] ^ m[90] ^ m[91] ^ m[92] ^ m[93] ^ m[94] ^ m[95] ^ m[96] ^ m[97] ^ m[98] ^ m[99] ^ m[100] ^ m[101] ^ m[102] ^ m[103] ^ m[104] ^ m[105] ^ m[106] ^ m[107] ^ m[108] ^ m[109] ^ m[110] ^ m[111] ^ m[112] ^ m[113] ^ m[114] ^ m[115] ^ m[116] ^ m[117] ^ m[118] ^ m[119] ^ m[156] ^ m[157] ^ m[158] ^ m[159] ^ m[160] ^ m[161] ^ m[162] ^ m[163] ^ m[164] ^ m[201] ^ m[202] ^ m[203] ^ m[204] ^ m[205] ^ m[206] ^ m[207] ^ m[208] ^ m[209] ^ m[219] ^ m[346] ^ m[347] ^ m[348] ^ m[349] ^ m[350] ^ m[351] ^ m[352] ^ m[353] ^ m[354] ^ m[355] ^ m[356] ^ m[357] ^ m[358] ^ m[359] ^ m[360] ^ m[361] ^ m[362] ^ m[363] ^ m[364] ^ m[365] ^ m[366] ^ m[367] ^ m[368] ^ m[369] ^ m[370] ^ m[371] ^ m[372] ^ m[373] ^ m[374] ^ m[375] ^ m[376] ^ m[377] ^ m[378] ^ m[379] ^ m[380] ^ m[381] ^ m[382] ^ m[383] ^ m[384] ^ m[385] ^ m[386] ^ m[387] ^ m[388] ^ m[389] ^ m[390] ^ m[391] ^ m[392] ^ m[393] ^ m[394] ^ m[395] ^ m[396] ^ m[397] ^ m[398] ^ m[399] ^ m[400] ^ m[401] ^ m[402] ^ m[403] ^ m[404] ^ m[405] ^ m[406] ^ m[407] ^ m[408] ^ m[409] ^ m[410] ^ m[411] ^ m[412] ^ m[413] ^ m[414] ^ m[415] ^ m[416] ^ m[417] ^ m[418] ^ m[419] ^ m[420] ^ m[421] ^ m[422] ^ m[423] ^ m[424] ^ m[425] ^ m[426] ^ m[427] ^ m[428] ^ m[429] ^ m[430] ^ m[431] ^ m[432] ^ m[433] ^ m[434] ^ m[435] ^ m[436] ^ m[437] ^ m[438] ^ m[439] ^ m[440] ^ m[441] ^ m[442] ^ m[443] ^ m[444] ^ m[445] ^ m[446] ^ m[447] ^ m[448] ^ m[449] ^ m[450] ^ m[451] ^ m[452] ^ m[453] ^ m[454] ^ m[455] ^ m[456] ^ m[457] ^ m[458] ^ m[459] ^ m[460] ^ m[461] ^ m[462] ^ m[463] ^ m[464] ^ m[465] ^ m[466] ^ m[467] ^ m[468] ^ m[469] ^ m[470] ^ m[471] ^ m[598] ^ m[599] ^ m[600] ^ m[601] ^ m[602] ^ m[603] ^ m[604] ^ m[605] ^ m[606] ^ m[607] ^ m[608] ^ m[609] ^ m[610] ^ m[611] ^ m[612] ^ m[613] ^ m[614] ^ m[615] ^ m[616] ^ m[617] ^ m[618] ^ m[619] ^ m[620] ^ m[621] ^ m[622] ^ m[623] ^ m[624] ^ m[625] ^ m[626] ^ m[627] ^ m[628] ^ m[629] ^ m[630] ^ m[631] ^ m[632] ^ m[633] ^ m[634] ^ m[635] ^ m[636] ^ m[637] ^ m[638] ^ m[639] ^ m[640] ^ m[641] ^ m[642] ^ m[643] ^ m[644] ^ m[645] ^ m[646] ^ m[647] ^ m[648] ^ m[649] ^ m[650] ^ m[651] ^ m[652] ^ m[653] ^ m[654] ^ m[655] ^ m[656] ^ m[657] ^ m[658] ^ m[659] ^ m[660] ^ m[661] ^ m[662] ^ m[663] ^ m[664] ^ m[665] ^ m[666] ^ m[667] ^ m[668] ^ m[669] ^ m[670] ^ m[671] ^ m[672] ^ m[673] ^ m[674] ^ m[675] ^ m[676] ^ m[677] ^ m[678] ^ m[679] ^ m[680] ^ m[681] ^ m[808] ^ m[809] ^ m[810] ^ m[811] ^ m[812] ^ m[813] ^ m[814] ^ m[815] ^ m[816] ^ m[817] ^ m[818] ^ m[819] ^ m[820] ^ m[821] ^ m[822] ^ m[823] ^ m[824] ^ m[825] ^ m[826] ^ m[827] ^ m[828] ^ m[829] ^ m[830] ^ m[831] ^ m[832] ^ m[833] ^ m[834] ^ m[835] ^ m[836] ^ m[837] ^ m[838] ^ m[839] ^ m[840] ^ m[841] ^ m[842] ^ m[843] ^ m[844] ^ m[845] ^ m[846] ^ m[847] ^ m[848] ^ m[849] ^ m[850] ^ m[851] ^ m[852] ^ m[853] ^ m[854] ^ m[855] ^ m[856] ^ m[857] ^ m[858] ^ m[859] ^ m[860] ^ m[861] ^ m[862] ^ m[863] ^ m[864] ^ m[865] ^ m[866] ^ m[867] ^ m[868] ^ m[869] ^ m[870] ^ m[871] ^ m[872] ^ m[873] ^ m[874] ^ m[875] ^ m[876] ^ m[877] ^ m[878] ^ m[879] ^ m[880] ^ m[881] ^ m[882] ^ m[883] ^ m[884] ^ m[885] ^ m[886] ^ m[887] ^ m[888] ^ m[889] ^ m[890] ^ m[891] ^ m[976] ^ m[977] ^ m[978] ^ m[979] ^ m[980] ^ m[981] ^ m[982] ^ m[983] ^ m[984] ^ m[985] ^ m[986] ^ m[987] ^ m[988] ^ m[989] ^ m[990] ^ m[991] ^ m[992] ^ m[993] ^ m[994] ^ m[995] ^ m[996] ^ m[997] ^ m[998] ^ m[999] ^ m[1000] ^ m[1001] ^ m[1002] ^ m[1003] ^ m[1004] ^ m[1005] ^ m[1006] ^ m[1007] ^ m[1008] ^ m[1009] ^ m[1010] ^ m[1011];
    assign parity[3] = m[56] ^ m[57] ^ m[58] ^ m[59] ^ m[60] ^ m[61] ^ m[62] ^ m[63] ^ m[64] ^ m[65] ^ m[66] ^ m[67] ^ m[68] ^ m[69] ^ m[70] ^ m[71] ^ m[72] ^ m[73] ^ m[74] ^ m[75] ^ m[76] ^ m[77] ^ m[78] ^ m[79] ^ m[80] ^ m[81] ^ m[82] ^ m[83] ^ m[112] ^ m[113] ^ m[114] ^ m[115] ^ m[116] ^ m[117] ^ m[118] ^ m[119] ^ m[148] ^ m[149] ^ m[150] ^ m[151] ^ m[152] ^ m[153] ^ m[154] ^ m[155] ^ m[164] ^ m[193] ^ m[194] ^ m[195] ^ m[196] ^ m[197] ^ m[198] ^ m[199] ^ m[200] ^ m[209] ^ m[218] ^ m[276] ^ m[277] ^ m[278] ^ m[279] ^ m[280] ^ m[281] ^ m[282] ^ m[283] ^ m[284] ^ m[285] ^ m[286] ^ m[287] ^ m[288] ^ m[289] ^ m[290] ^ m[291] ^ m[292] ^ m[293] ^ m[294] ^ m[295] ^ m[296] ^ m[297] ^ m[298] ^ m[299] ^ m[300] ^ m[301] ^ m[302] ^ m[303] ^ m[304] ^ m[305] ^ m[306] ^ m[307] ^ m[308] ^ m[309] ^ m[310] ^ m[311] ^ m[312] ^ m[313] ^ m[314] ^ m[315] ^ m[316] ^ m[317] ^ m[318] ^ m[319] ^ m[320] ^ m[321] ^ m[322] ^ m[323] ^ m[324] ^ m[325] ^ m[326] ^ m[327] ^ m[328] ^ m[329] ^ m[330] ^ m[331] ^ m[332] ^ m[333] ^ m[334] ^ m[335] ^ m[336] ^ m[337] ^ m[338] ^ m[339] ^ m[340] ^ m[341] ^ m[342] ^ m[343] ^ m[344] ^ m[345] ^ m[416] ^ m[417] ^ m[418] ^ m[419] ^ m[420] ^ m[421] ^ m[422] ^ m[423] ^ m[424] ^ m[425] ^ m[426] ^ m[427] ^ m[428] ^ m[429] ^ m[430] ^ m[431] ^ m[432] ^ m[433] ^ m[434] ^ m[435] ^ m[436] ^ m[437] ^ m[438] ^ m[439] ^ m[440] ^ m[441] ^ m[442] ^ m[443] ^ m[444] ^ m[445] ^ m[446] ^ m[447] ^ m[448] ^ m[449] ^ m[450] ^ m[451] ^ m[452] ^ m[453] ^ m[454] ^ m[455] ^ m[456] ^ m[457] ^ m[458] ^ m[459] ^ m[460] ^ m[461] ^ m[462] ^ m[463] ^ m[464] ^ m[465] ^ m[466] ^ m[467] ^ m[468] ^ m[469] ^ m[470] ^ m[471] ^ m[542] ^ m[543] ^ m[544] ^ m[545] ^ m[546] ^ m[547] ^ m[548] ^ m[549] ^ m[550] ^ m[551] ^ m[552] ^ m[553] ^ m[554] ^ m[555] ^ m[556] ^ m[557] ^ m[558] ^ m[559] ^ m[560] ^ m[561] ^ m[562] ^ m[563] ^ m[564] ^ m[565] ^ m[566] ^ m[567] ^ m[568] ^ m[569] ^ m[570] ^ m[571] ^ m[572] ^ m[573] ^ m[574] ^ m[575] ^ m[576] ^ m[577] ^ m[578] ^ m[579] ^ m[580] ^ m[581] ^ m[582] ^ m[583] ^ m[584] ^ m[585] ^ m[586] ^ m[587] ^ m[588] ^ m[589] ^ m[590] ^ m[591] ^ m[592] ^ m[593] ^ m[594] ^ m[595] ^ m[596] ^ m[597] ^ m[654] ^ m[655] ^ m[656] ^ m[657] ^ m[658] ^ m[659] ^ m[660] ^ m[661] ^ m[662] ^ m[663] ^ m[664] ^ m[665] ^ m[666] ^ m[667] ^ m[668] ^ m[669] ^ m[670] ^ m[671] ^ m[672] ^ m[673] ^ m[674] ^ m[675] ^ m[676] ^ m[677] ^ m[678] ^ m[679] ^ m[680] ^ m[681] ^ m[752] ^ m[753] ^ m[754] ^ m[755] ^ m[756] ^ m[757] ^ m[758] ^ m[759] ^ m[760] ^ m[761] ^ m[762] ^ m[763] ^ m[764] ^ m[765] ^ m[766] ^ m[767] ^ m[768] ^ m[769] ^ m[770] ^ m[771] ^ m[772] ^ m[773] ^ m[774] ^ m[775] ^ m[776] ^ m[777] ^ m[778] ^ m[779] ^ m[780] ^ m[781] ^ m[782] ^ m[783] ^ m[784] ^ m[785] ^ m[786] ^ m[787] ^ m[788] ^ m[789] ^ m[790] ^ m[791] ^ m[792] ^ m[793] ^ m[794] ^ m[795] ^ m[796] ^ m[797] ^ m[798] ^ m[799] ^ m[800] ^ m[801] ^ m[802] ^ m[803] ^ m[804] ^ m[805] ^ m[806] ^ m[807] ^ m[864] ^ m[865] ^ m[866] ^ m[867] ^ m[868] ^ m[869] ^ m[870] ^ m[871] ^ m[872] ^ m[873] ^ m[874] ^ m[875] ^ m[876] ^ m[877] ^ m[878] ^ m[879] ^ m[880] ^ m[881] ^ m[882] ^ m[883] ^ m[884] ^ m[885] ^ m[886] ^ m[887] ^ m[888] ^ m[889] ^ m[890] ^ m[891] ^ m[948] ^ m[949] ^ m[950] ^ m[951] ^ m[952] ^ m[953] ^ m[954] ^ m[955] ^ m[956] ^ m[957] ^ m[958] ^ m[959] ^ m[960] ^ m[961] ^ m[962] ^ m[963] ^ m[964] ^ m[965] ^ m[966] ^ m[967] ^ m[968] ^ m[969] ^ m[970] ^ m[971] ^ m[972] ^ m[973] ^ m[974] ^ m[975] ^ m[1004] ^ m[1005] ^ m[1006] ^ m[1007] ^ m[1008] ^ m[1009] ^ m[1010] ^ m[1011] ^ m[1020] ^ m[1021] ^ m[1022] ^ m[1023];
    assign parity[4] = m[35] ^ m[36] ^ m[37] ^ m[38] ^ m[39] ^ m[40] ^ m[41] ^ m[42] ^ m[43] ^ m[44] ^ m[45] ^ m[46] ^ m[47] ^ m[48] ^ m[49] ^ m[50] ^ m[51] ^ m[52] ^ m[53] ^ m[54] ^ m[55] ^ m[77] ^ m[78] ^ m[79] ^ m[80] ^ m[81] ^ m[82] ^ m[83] ^ m[105] ^ m[106] ^ m[107] ^ m[108] ^ m[109] ^ m[110] ^ m[111] ^ m[119] ^ m[141] ^ m[142] ^ m[143] ^ m[144] ^ m[145] ^ m[146] ^ m[147] ^ m[155] ^ m[163] ^ m[186] ^ m[187] ^ m[188] ^ m[189] ^ m[190] ^ m[191] ^ m[192] ^ m[200] ^ m[208] ^ m[217] ^ m[241] ^ m[242] ^ m[243] ^ m[244] ^ m[245] ^ m[246] ^ m[247] ^ m[248] ^ m[249] ^ m[250] ^ m[251] ^ m[252] ^ m[253] ^ m[254] ^ m[255] ^ m[256] ^ m[257] ^ m[258] ^ m[259] ^ m[260] ^ m[261] ^ m[262] ^ m[263] ^ m[264] ^ m[265] ^ m[266] ^ m[267] ^ m[268] ^ m[269] ^ m[270] ^ m[271] ^ m[272] ^ m[273] ^ m[274] ^ m[275] ^ m[311] ^ m[312] ^ m[313] ^ m[314] ^ m[315] ^ m[316] ^ m[317] ^ m[318] ^ m[319] ^ m[320] ^ m[321] ^ m[322] ^ m[323] ^ m[324] ^ m[325] ^ m[326] ^ m[327] ^ m[328] ^ m[329] ^ m[330] ^ m[331] ^ m[332] ^ m[333] ^ m[334] ^ m[335] ^ m[336] ^ m[337] ^ m[338] ^ m[339] ^ m[340] ^ m[341] ^ m[342] ^ m[343] ^ m[344] ^ m[345] ^ m[381] ^ m[382] ^ m[383] ^ m[384] ^ m[385] ^ m[386] ^ m[387] ^ m[388] ^ m[389] ^ m[390] ^ m[391] ^ m[392] ^ m[393] ^ m[394] ^ m[395] ^ m[396] ^ m[397] ^ m[398] ^ m[399] ^ m[400] ^ m[401] ^ m[402] ^ m[403] ^ m[404] ^ m[405] ^ m[406] ^ m[407] ^ m[408] ^ m[409] ^ m[410] ^ m[411] ^ m[412] ^ m[413] ^ m[414] ^ m[415] ^ m[451] ^ m[452] ^ m[453] ^ m[454] ^ m[455] ^ m[456] ^ m[457] ^ m[458] ^ m[459] ^ m[460] ^ m[461] ^ m[462] ^ m[463] ^ m[464] ^ m[465] ^ m[466] ^ m[467] ^ m[468] ^ m[469] ^ m[470] ^ m[471] ^ m[507] ^ m[508] ^ m[509] ^ m[510] ^ m[511] ^ m[512] ^ m[513] ^ m[514] ^ m[515] ^ m[516] ^ m[517] ^ m[518] ^ m[519] ^ m[520] ^ m[521] ^ m[522] ^ m[523] ^ m[524] ^ m[525] ^ m[526] ^ m[527] ^ m[528] ^ m[529] ^ m[530] ^ m[531] ^ m[532] ^ m[533] ^ m[534] ^ m[535] ^ m[536] ^ m[537] ^ m[538] ^ m[539] ^ m[540] ^ m[541] ^ m[577] ^ m[578] ^ m[579] ^ m[580] ^ m[581] ^ m[582] ^ m[583] ^ m[584] ^ m[585] ^ m[586] ^ m[587] ^ m[588] ^ m[589] ^ m[590] ^ m[591] ^ m[592] ^ m[593] ^ m[594] ^ m[595] ^ m[596] ^ m[597] ^ m[633] ^ m[634] ^ m[635] ^ m[636] ^ m[637] ^ m[638] ^ m[639] ^ m[640] ^ m[641] ^ m[642] ^ m[643] ^ m[644] ^ m[645] ^ m[646] ^ m[647] ^ m[648] ^ m[649] ^ m[650] ^ m[651] ^ m[652] ^ m[653] ^ m[675] ^ m[676] ^ m[677] ^ m[678] ^ m[679] ^ m[680] ^ m[681] ^ m[717] ^ m[718] ^ m[719] ^ m[720] ^ m[721] ^ m[722] ^ m[723] ^ m[724] ^ m[725] ^ m[726] ^ m[727] ^ m[728] ^ m[729] ^ m[730] ^ m[731] ^ m[732] ^ m[733] ^ m[734] ^ m[735] ^ m[736] ^ m[737] ^ m[738] ^ m[739] ^ m[740] ^ m[741] ^ m[742] ^ m[743] ^ m[744] ^ m[745] ^ m[746] ^ m[747] ^ m[748] ^ m[749] ^ m[750] ^ m[751] ^ m[787] ^ m[788] ^ m[789] ^ m[790] ^ m[791] ^ m[792] ^ m[793] ^ m[794] ^ m[795] ^ m[796] ^ m[797] ^ m[798] ^ m[799] ^ m[800] ^ m[801] ^ m[802] ^ m[803] ^ m[804] ^ m[805] ^ m[806] ^ m[807] ^ m[843] ^ m[844] ^ m[845] ^ m[846] ^ m[847] ^ m[848] ^ m[849] ^ m[850] ^ m[851] ^ m[852] ^ m[853] ^ m[854] ^ m[855] ^ m[856] ^ m[857] ^ m[858] ^ m[859] ^ m[860] ^ m[861] ^ m[862] ^ m[863] ^ m[885] ^ m[886] ^ m[887] ^ m[888] ^ m[889] ^ m[890] ^ m[891] ^ m[927] ^ m[928] ^ m[929] ^ m[930] ^ m[931] ^ m[932] ^ m[933] ^ m[934] ^ m[935] ^ m[936] ^ m[937] ^ m[938] ^ m[939] ^ m[940] ^ m[941] ^ m[942] ^ m[943] ^ m[944] ^ m[945] ^ m[946] ^ m[947] ^ m[969] ^ m[970] ^ m[971] ^ m[972] ^ m[973] ^ m[974] ^ m[975] ^ m[997] ^ m[998] ^ m[999] ^ m[1000] ^ m[1001] ^ m[1002] ^ m[1003] ^ m[1011] ^ m[1013] ^ m[1014] ^ m[1015] ^ m[1016] ^ m[1017] ^ m[1018] ^ m[1019];
    assign parity[5] = m[20] ^ m[21] ^ m[22] ^ m[23] ^ m[24] ^ m[25] ^ m[26] ^ m[27] ^ m[28] ^ m[29] ^ m[30] ^ m[31] ^ m[32] ^ m[33] ^ m[34] ^ m[50] ^ m[51] ^ m[52] ^ m[53] ^ m[54] ^ m[55] ^ m[71] ^ m[72] ^ m[73] ^ m[74] ^ m[75] ^ m[76] ^ m[83] ^ m[99] ^ m[100] ^ m[101] ^ m[102] ^ m[103] ^ m[104] ^ m[111] ^ m[118] ^ m[135] ^ m[136] ^ m[137] ^ m[138] ^ m[139] ^ m[140] ^ m[147] ^ m[154] ^ m[162] ^ m[180] ^ m[181] ^ m[182] ^ m[183] ^ m[184] ^ m[185] ^ m[192] ^ m[199] ^ m[207] ^ m[216] ^ m[226] ^ m[227] ^ m[228] ^ m[229] ^ m[230] ^ m[231] ^ m[232] ^ m[233] ^ m[234] ^ m[235] ^ m[236] ^ m[237] ^ m[238] ^ m[239] ^ m[240] ^ m[256] ^ m[257] ^ m[258] ^ m[259] ^ m[260] ^ m[261] ^ m[262] ^ m[263] ^ m[264] ^ m[265] ^ m[266] ^ m[267] ^ m[268] ^ m[269] ^ m[270] ^ m[271] ^ m[272] ^ m[273] ^ m[274] ^ m[275] ^ m[291] ^ m[292] ^ m[293] ^ m[294] ^ m[295] ^ m[296] ^ m[297] ^ m[298] ^ m[299] ^ m[300] ^ m[301] ^ m[302] ^ m[303] ^ m[304] ^ m[305] ^ m[306] ^ m[307] ^ m[308] ^ m[309] ^ m[310] ^ m[331] ^ m[332] ^ m[333] ^ m[334] ^ m[335] ^ m[336] ^ m[337] ^ m[338] ^ m[339] ^ m[340] ^ m[341] ^ m[342] ^ m[343] ^ m[344] ^ m[345] ^ m[361] ^ m[362] ^ m[363] ^ m[364] ^ m[365] ^ m[366] ^ m[367] ^ m[368] ^ m[369] ^ m[370] ^ m[371] ^ m[372] ^ m[373] ^ m[374] ^ m[375] ^ m[376] ^ m[377] ^ m[378] ^ m[379] ^ m[380] ^ m[401] ^ m[402] ^ m[403] ^ m[404] ^ m[405] ^ m[406] ^ m[407] ^ m[408] ^ m[409] ^ m[410] ^ m[411] ^ m[412] ^ m[413] ^ m[414] ^ m[415] ^ m[436] ^ m[437] ^ m[438] ^ m[439] ^ m[440] ^ m[441] ^ m[442] ^ m[443] ^ m[444] ^ m[445] ^ m[446] ^ m[447] ^ m[448] ^ m[449] ^ m[450] ^ m[466] ^ m[467] ^ m[468] ^ m[469] ^ m[470] ^ m[471] ^ m[487] ^ m[488] ^ m[489] ^ m[490] ^ m[491] ^ m[492] ^ m[493] ^ m[494] ^ m[495] ^ m[496] ^ m[497] ^ m[498] ^ m[499] ^ m[500] ^ m[501] ^ m[502] ^ m[503] ^ m[504] ^ m[505] ^ m[506] ^ m[527] ^ m[528] ^ m[529] ^ m[530] ^ m[531] ^ m[532] ^ m[533] ^ m[534] ^ m[535] ^ m[536] ^ m[537] ^ m[538] ^ m[539] ^ m[540] ^ m[541] ^ m[562] ^ m[563] ^ m[564] ^ m[565] ^ m[566] ^ m[567] ^ m[568] ^ m[569] ^ m[570] ^ m[571] ^ m[572] ^ m[573] ^ m[574] ^ m[575] ^ m[576] ^ m[592] ^ m[593] ^ m[594] ^ m[595] ^ m[596] ^ m[597] ^ m[618] ^ m[619] ^ m[620] ^ m[621] ^ m[622] ^ m[623] ^ m[624] ^ m[625] ^ m[626] ^ m[627] ^ m[628] ^ m[629] ^ m[630] ^ m[631] ^ m[632] ^ m[648] ^ m[649] ^ m[650] ^ m[651] ^ m[652] ^ m[653] ^ m[669] ^ m[670] ^ m[671] ^ m[672] ^ m[673] ^ m[674] ^ m[681] ^ m[697] ^ m[698] ^ m[699] ^ m[700] ^ m[701] ^ m[702] ^ m[703] ^ m[704] ^ m[705] ^ m[706] ^ m[707] ^ m[708] ^ m[709] ^ m[710] ^ m[711] ^ m[712] ^ m[713] ^ m[714] ^ m[715] ^ m[716] ^ m[737] ^ m[738] ^ m[739] ^ m[740] ^ m[741] ^ m[742] ^ m[743] ^ m[744] ^ m[745] ^ m[746] ^ m[747] ^ m[748] ^ m[749] ^ m[750] ^ m[751] ^ m[772] ^ m[773] ^ m[774] ^ m[775] ^ m[776] ^ m[777] ^ m[778] ^ m[779] ^ m[780] ^ m[781] ^ m[782] ^ m[783] ^ m[784] ^ m[785] ^ m[786] ^ m[802] ^ m[803] ^ m[804] ^ m[805] ^ m[806] ^ m[807] ^ m[828] ^ m[829] ^ m[830] ^ m[831] ^ m[832] ^ m[833] ^ m[834] ^ m[835] ^ m[836] ^ m[837] ^ m[838] ^ m[839] ^ m[840] ^ m[841] ^ m[842] ^ m[858] ^ m[859] ^ m[860] ^ m[861] ^ m[862] ^ m[863] ^ m[879] ^ m[880] ^ m[881] ^ m[882] ^ m[883] ^ m[884] ^ m[891] ^ m[912] ^ m[913] ^ m[914] ^ m[915] ^ m[916] ^ m[917] ^ m[918] ^ m[919] ^ m[920] ^ m[921] ^ m[922] ^ m[923] ^ m[924] ^ m[925] ^ m[926] ^ m[942] ^ m[943] ^ m[944] ^ m[945] ^ m[946] ^ m[947] ^ m[963] ^ m[964] ^ m[965] ^ m[966] ^ m[967] ^ m[968] ^ m[975] ^ m[991] ^ m[992] ^ m[993] ^ m[994] ^ m[995] ^ m[996] ^ m[1003] ^ m[1010] ^ m[1012] ^ m[1014] ^ m[1015] ^ m[1016] ^ m[1017] ^ m[1018] ^ m[1019] ^ m[1021] ^ m[1022] ^ m[1023];
    assign parity[6] = m[10] ^ m[11] ^ m[12] ^ m[13] ^ m[14] ^ m[15] ^ m[16] ^ m[17] ^ m[18] ^ m[19] ^ m[30] ^ m[31] ^ m[32] ^ m[33] ^ m[34] ^ m[45] ^ m[46] ^ m[47] ^ m[48] ^ m[49] ^ m[55] ^ m[66] ^ m[67] ^ m[68] ^ m[69] ^ m[70] ^ m[76] ^ m[82] ^ m[94] ^ m[95] ^ m[96] ^ m[97] ^ m[98] ^ m[104] ^ m[110] ^ m[117] ^ m[130] ^ m[131] ^ m[132] ^ m[133] ^ m[134] ^ m[140] ^ m[146] ^ m[153] ^ m[161] ^ m[175] ^ m[176] ^ m[177] ^ m[178] ^ m[179] ^ m[185] ^ m[191] ^ m[198] ^ m[206] ^ m[215] ^ m[221] ^ m[222] ^ m[223] ^ m[224] ^ m[225] ^ m[231] ^ m[232] ^ m[233] ^ m[234] ^ m[235] ^ m[236] ^ m[237] ^ m[238] ^ m[239] ^ m[240] ^ m[246] ^ m[247] ^ m[248] ^ m[249] ^ m[250] ^ m[251] ^ m[252] ^ m[253] ^ m[254] ^ m[255] ^ m[266] ^ m[267] ^ m[268] ^ m[269] ^ m[270] ^ m[271] ^ m[272] ^ m[273] ^ m[274] ^ m[275] ^ m[281] ^ m[282] ^ m[283] ^ m[284] ^ m[285] ^ m[286] ^ m[287] ^ m[288] ^ m[289] ^ m[290] ^ m[301] ^ m[302] ^ m[303] ^ m[304] ^ m[305] ^ m[306] ^ m[307] ^ m[308] ^ m[309] ^ m[310] ^ m[321] ^ m[322] ^ m[323] ^ m[324] ^ m[325] ^ m[326] ^ m[327] ^ m[328] ^ m[329] ^ m[330] ^ m[341] ^ m[342] ^ m[343] ^ m[344] ^ m[345] ^ m[351] ^ m[352] ^ m[353] ^ m[354] ^ m[355] ^ m[356] ^ m[357] ^ m[358] ^ m[359] ^ m[360] ^ m[371] ^ m[372] ^ m[373] ^ m[374] ^ m[375] ^ m[376] ^ m[377] ^ m[378] ^ m[379] ^ m[380] ^ m[391] ^ m[392] ^ m[393] ^ m[394] ^ m[395] ^ m[396] ^ m[397] ^ m[398] ^ m[399] ^ m[400] ^ m[411] ^ m[412] ^ m[413] ^ m[414] ^ m[415] ^ m[426] ^ m[427] ^ m[428] ^ m[429] ^ m[430] ^ m[431] ^ m[432] ^ m[433] ^ m[434] ^ m[435] ^ m[446] ^ m[447] ^ m[448] ^ m[449] ^ m[450] ^ m[461] ^ m[462] ^ m[463] ^ m[464] ^ m[465] ^ m[471] ^ m[477] ^ m[478] ^ m[479] ^ m[480] ^ m[481] ^ m[482] ^ m[483] ^ m[484] ^ m[485] ^ m[486] ^ m[497] ^ m[498] ^ m[499] ^ m[500] ^ m[501] ^ m[502] ^ m[503] ^ m[504] ^ m[505] ^ m[506] ^ m[517] ^ m[518] ^ m[519] ^ m[520] ^ m[521] ^ m[522] ^ m[523] ^ m[524] ^ m[525] ^ m[526] ^ m[537] ^ m[538] ^ m[539] ^ m[540] ^ m[541] ^ m[552] ^ m[553] ^ m[554] ^ m[555] ^ m[556] ^ m[557] ^ m[558] ^ m[559] ^ m[560] ^ m[561] ^ m[572] ^ m[573] ^ m[574] ^ m[575] ^ m[576] ^ m[587] ^ m[588] ^ m[589] ^ m[590] ^ m[591] ^ m[597] ^ m[608] ^ m[609] ^ m[610] ^ m[611] ^ m[612] ^ m[613] ^ m[614] ^ m[615] ^ m[616] ^ m[617] ^ m[628] ^ m[629] ^ m[630] ^ m[631] ^ m[632] ^ m[643] ^ m[644] ^ m[645] ^ m[646] ^ m[647] ^ m[653] ^ m[664] ^ m[665] ^ m[666] ^ m[667] ^ m[668] ^ m[674] ^ m[680] ^ m[687] ^ m[688] ^ m[689] ^ m[690] ^ m[691] ^ m[692] ^ m[693] ^ m[694] ^ m[695] ^ m[696] ^ m[707] ^ m[708] ^ m[709] ^ m[710] ^ m[711] ^ m[712] ^ m[713] ^ m[714] ^ m[715] ^ m[716] ^ m[727] ^ m[728] ^ m[729] ^ m[730] ^ m[731] ^ m[732] ^ m[733] ^ m[734] ^ m[735] ^ m[736] ^ m[747] ^ m[748] ^ m[749] ^ m[750] ^ m[751] ^ m[762] ^ m[763] ^ m[764] ^ m[765] ^ m[766] ^ m[767] ^ m[768] ^ m[769] ^ m[770] ^ m[771] ^ m[782] ^ m[783] ^ m[784] ^ m[785] ^ m[786] ^ m[797] ^ m[798] ^ m[799] ^ m[800] ^ m[801] ^ m[807] ^ m[818] ^ m[819] ^ m[820] ^ m[821] ^ m[822] ^ m[823] ^ m[824] ^ m[825] ^ m[826] ^ m[827] ^ m[838] ^ m[839] ^ m[840] ^ m[841] ^ m[842] ^ m[853] ^ m[854] ^ m[855] ^ m[856] ^ m[857] ^ m[863] ^ m[874] ^ m[875] ^ m[876] ^ m[877] ^ m[878] ^ m[884] ^ m[890] ^ m[902] ^ m[903] ^ m[904] ^ m[905] ^ m[906] ^ m[907] ^ m[908] ^ m[909] ^ m[910] ^ m[911] ^ m[922] ^ m[923] ^ m[924] ^ m[925] ^ m[926] ^ m[937] ^ m[938] ^ m[939] ^ m[940] ^ m[941] ^ m[947] ^ m[958] ^ m[959] ^ m[960] ^ m[961] ^ m[962] ^ m[968] ^ m[974] ^ m[986] ^ m[987] ^ m[988] ^ m[989] ^ m[990] ^ m[996] ^ m[1002] ^ m[1009] ^ m[1012] ^ m[1013] ^ m[1015] ^ m[1016] ^ m[1017] ^ m[1018] ^ m[1019] ^ m[1020] ^ m[1022] ^ m[1023];
    assign parity[7] = m[4] ^ m[5] ^ m[6] ^ m[7] ^ m[8] ^ m[9] ^ m[16] ^ m[17] ^ m[18] ^ m[19] ^ m[26] ^ m[27] ^ m[28] ^ m[29] ^ m[34] ^ m[41] ^ m[42] ^ m[43] ^ m[44] ^ m[49] ^ m[54] ^ m[62] ^ m[63] ^ m[64] ^ m[65] ^ m[70] ^ m[75] ^ m[81] ^ m[90] ^ m[91] ^ m[92] ^ m[93] ^ m[98] ^ m[103] ^ m[109] ^ m[116] ^ m[126] ^ m[127] ^ m[128] ^ m[129] ^ m[134] ^ m[139] ^ m[145] ^ m[152] ^ m[160] ^ m[171] ^ m[172] ^ m[173] ^ m[174] ^ m[179] ^ m[184] ^ m[190] ^ m[197] ^ m[205] ^ m[214] ^ m[220] ^ m[222] ^ m[223] ^ m[224] ^ m[225] ^ m[227] ^ m[228] ^ m[229] ^ m[230] ^ m[235] ^ m[236] ^ m[237] ^ m[238] ^ m[239] ^ m[240] ^ m[242] ^ m[243] ^ m[244] ^ m[245] ^ m[250] ^ m[251] ^ m[252] ^ m[253] ^ m[254] ^ m[255] ^ m[260] ^ m[261] ^ m[262] ^ m[263] ^ m[264] ^ m[265] ^ m[272] ^ m[273] ^ m[274] ^ m[275] ^ m[277] ^ m[278] ^ m[279] ^ m[280] ^ m[285] ^ m[286] ^ m[287] ^ m[288] ^ m[289] ^ m[290] ^ m[295] ^ m[296] ^ m[297] ^ m[298] ^ m[299] ^ m[300] ^ m[307] ^ m[308] ^ m[309] ^ m[310] ^ m[315] ^ m[316] ^ m[317] ^ m[318] ^ m[319] ^ m[320] ^ m[327] ^ m[328] ^ m[329] ^ m[330] ^ m[337] ^ m[338] ^ m[339] ^ m[340] ^ m[345] ^ m[347] ^ m[348] ^ m[349] ^ m[350] ^ m[355] ^ m[356] ^ m[357] ^ m[358] ^ m[359] ^ m[360] ^ m[365] ^ m[366] ^ m[367] ^ m[368] ^ m[369] ^ m[370] ^ m[377] ^ m[378] ^ m[379] ^ m[380] ^ m[385] ^ m[386] ^ m[387] ^ m[388] ^ m[389] ^ m[390] ^ m[397] ^ m[398] ^ m[399] ^ m[400] ^ m[407] ^ m[408] ^ m[409] ^ m[410] ^ m[415] ^ m[420] ^ m[421] ^ m[422] ^ m[423] ^ m[424] ^ m[425] ^ m[432] ^ m[433] ^ m[434] ^ m[435] ^ m[442] ^ m[443] ^ m[444] ^ m[445] ^ m[450] ^ m[457] ^ m[458] ^ m[459] ^ m[460] ^ m[465] ^ m[470] ^ m[473] ^ m[474] ^ m[475] ^ m[476] ^ m[481] ^ m[482] ^ m[483] ^ m[484] ^ m[485] ^ m[486] ^ m[491] ^ m[492] ^ m[493] ^ m[494] ^ m[495] ^ m[496] ^ m[503] ^ m[504] ^ m[505] ^ m[506] ^ m[511] ^ m[512] ^ m[513] ^ m[514] ^ m[515] ^ m[516] ^ m[523] ^ m[524] ^ m[525] ^ m[526] ^ m[533] ^ m[534] ^ m[535] ^ m[536] ^ m[541] ^ m[546] ^ m[547] ^ m[548] ^ m[549] ^ m[550] ^ m[551] ^ m[558] ^ m[559] ^ m[560] ^ m[561] ^ m[568] ^ m[569] ^ m[570] ^ m[571] ^ m[576] ^ m[583] ^ m[584] ^ m[585] ^ m[586] ^ m[591] ^ m[596] ^ m[602] ^ m[603] ^ m[604] ^ m[605] ^ m[606] ^ m[607] ^ m[614] ^ m[615] ^ m[616] ^ m[617] ^ m[624] ^ m[625] ^ m[626] ^ m[627] ^ m[632] ^ m[639] ^ m[640] ^ m[641] ^ m[642] ^ m[647] ^ m[652] ^ m[660] ^ m[661] ^ m[662] ^ m[663] ^ m[668] ^ m[673] ^ m[679] ^ m[683] ^ m[684] ^ m[685] ^ m[686] ^ m[691] ^ m[692] ^ m[693] ^ m[694] ^ m[695] ^ m[696] ^ m[701] ^ m[702] ^ m[703] ^ m[704] ^ m[705] ^ m[706] ^ m[713] ^ m[714] ^ m[715] ^ m[716] ^ m[721] ^ m[722] ^ m[723] ^ m[724] ^ m[725] ^ m[726] ^ m[733] ^ m[734] ^ m[735] ^ m[736] ^ m[743] ^ m[744] ^ m[745] ^ m[746] ^ m[751] ^ m[756] ^ m[757] ^ m[758] ^ m[759] ^ m[760] ^ m[761] ^ m[768] ^ m[769] ^ m[770] ^ m[771] ^ m[778] ^ m[779] ^ m[780] ^ m[781] ^ m[786] ^ m[793] ^ m[794] ^ m[795] ^ m[796] ^ m[801] ^ m[806] ^ m[812] ^ m[813] ^ m[814] ^ m[815] ^ m[816] ^ m[817] ^ m[824] ^ m[825] ^ m[826] ^ m[827] ^ m[834] ^ m[835] ^ m[836] ^ m[837] ^ m[842] ^ m[849] ^ m[850] ^ m[851] ^ m[852] ^ m[857] ^ m[862] ^ m[870] ^ m[871] ^ m[872] ^ m[873] ^ m[878] ^ m[883] ^ m[889] ^ m[896] ^ m[897] ^ m[898] ^ m[899] ^ m[900] ^ m[901] ^ m[908] ^ m[909] ^ m[910] ^ m[911] ^ m[918] ^ m[919] ^ m[920] ^ m[921] ^ m[926] ^ m[933] ^ m[934] ^ m[935] ^ m[936] ^ m[941] ^ m[946] ^ m[954] ^ m[955] ^ m[956] ^ m[957] ^ m[962] ^ m[967] ^ m[973] ^ m[982] ^ m[983] ^ m[984] ^ m[985] ^ m[990] ^ m[995] ^ m[1001] ^ m[1008] ^ m[1012] ^ m[1013] ^ m[1014] ^ m[1016] ^ m[1017] ^ m[1018] ^ m[1019] ^ m[1020] ^ m[1021] ^ m[1023];
    assign parity[8] = m[1] ^ m[2] ^ m[3] ^ m[7] ^ m[8] ^ m[9] ^ m[13] ^ m[14] ^ m[15] ^ m[19] ^ m[23] ^ m[24] ^ m[25] ^ m[29] ^ m[33] ^ m[38] ^ m[39] ^ m[40] ^ m[44] ^ m[48] ^ m[53] ^ m[59] ^ m[60] ^ m[61] ^ m[65] ^ m[69] ^ m[74] ^ m[80] ^ m[87] ^ m[88] ^ m[89] ^ m[93] ^ m[97] ^ m[102] ^ m[108] ^ m[115] ^ m[123] ^ m[124] ^ m[125] ^ m[129] ^ m[133] ^ m[138] ^ m[144] ^ m[151] ^ m[159] ^ m[168] ^ m[169] ^ m[170] ^ m[174] ^ m[178] ^ m[183] ^ m[189] ^ m[196] ^ m[204] ^ m[213] ^ m[220] ^ m[221] ^ m[223] ^ m[224] ^ m[225] ^ m[226] ^ m[228] ^ m[229] ^ m[230] ^ m[232] ^ m[233] ^ m[234] ^ m[238] ^ m[239] ^ m[240] ^ m[241] ^ m[243] ^ m[244] ^ m[245] ^ m[247] ^ m[248] ^ m[249] ^ m[253] ^ m[254] ^ m[255] ^ m[257] ^ m[258] ^ m[259] ^ m[263] ^ m[264] ^ m[265] ^ m[269] ^ m[270] ^ m[271] ^ m[275] ^ m[276] ^ m[278] ^ m[279] ^ m[280] ^ m[282] ^ m[283] ^ m[284] ^ m[288] ^ m[289] ^ m[290] ^ m[292] ^ m[293] ^ m[294] ^ m[298] ^ m[299] ^ m[300] ^ m[304] ^ m[305] ^ m[306] ^ m[310] ^ m[312] ^ m[313] ^ m[314] ^ m[318] ^ m[319] ^ m[320] ^ m[324] ^ m[325] ^ m[326] ^ m[330] ^ m[334] ^ m[335] ^ m[336] ^ m[340] ^ m[344] ^ m[346] ^ m[348] ^ m[349] ^ m[350] ^ m[352] ^ m[353] ^ m[354] ^ m[358] ^ m[359] ^ m[360] ^ m[362] ^ m[363] ^ m[364] ^ m[368] ^ m[369] ^ m[370] ^ m[374] ^ m[375] ^ m[376] ^ m[380] ^ m[382] ^ m[383] ^ m[384] ^ m[388] ^ m[389] ^ m[390] ^ m[394] ^ m[395] ^ m[396] ^ m[400] ^ m[404] ^ m[405] ^ m[406] ^ m[410] ^ m[414] ^ m[417] ^ m[418] ^ m[419] ^ m[423] ^ m[424] ^ m[425] ^ m[429] ^ m[430] ^ m[431] ^ m[435] ^ m[439] ^ m[440] ^ m[441] ^ m[445] ^ m[449] ^ m[454] ^ m[455] ^ m[456] ^ m[460] ^ m[464] ^ m[469] ^ m[472] ^ m[474] ^ m[475] ^ m[476] ^ m[478] ^ m[479] ^ m[480] ^ m[484] ^ m[485] ^ m[486] ^ m[488] ^ m[489] ^ m[490] ^ m[494] ^ m[495] ^ m[496] ^ m[500] ^ m[501] ^ m[502] ^ m[506] ^ m[508] ^ m[509] ^ m[510] ^ m[514] ^ m[515] ^ m[516] ^ m[520] ^ m[521] ^ m[522] ^ m[526] ^ m[530] ^ m[531] ^ m[532] ^ m[536] ^ m[540] ^ m[543] ^ m[544] ^ m[545] ^ m[549] ^ m[550] ^ m[551] ^ m[555] ^ m[556] ^ m[557] ^ m[561] ^ m[565] ^ m[566] ^ m[567] ^ m[571] ^ m[575] ^ m[580] ^ m[581] ^ m[582] ^ m[586] ^ m[590] ^ m[595] ^ m[599] ^ m[600] ^ m[601] ^ m[605] ^ m[606] ^ m[607] ^ m[611] ^ m[612] ^ m[613] ^ m[617] ^ m[621] ^ m[622] ^ m[623] ^ m[627] ^ m[631] ^ m[636] ^ m[637] ^ m[638] ^ m[642] ^ m[646] ^ m[651] ^ m[657] ^ m[658] ^ m[659] ^ m[663] ^ m[667] ^ m[672] ^ m[678] ^ m[682] ^ m[684] ^ m[685] ^ m[686] ^ m[688] ^ m[689] ^ m[690] ^ m[694] ^ m[695] ^ m[696] ^ m[698] ^ m[699] ^ m[700] ^ m[704] ^ m[705] ^ m[706] ^ m[710] ^ m[711] ^ m[712] ^ m[716] ^ m[718] ^ m[719] ^ m[720] ^ m[724] ^ m[725] ^ m[726] ^ m[730] ^ m[731] ^ m[732] ^ m[736] ^ m[740] ^ m[741] ^ m[742] ^ m[746] ^ m[750] ^ m[753] ^ m[754] ^ m[755] ^ m[759] ^ m[760] ^ m[761] ^ m[765] ^ m[766] ^ m[767] ^ m[771] ^ m[775] ^ m[776] ^ m[777] ^ m[781] ^ m[785] ^ m[790] ^ m[791] ^ m[792] ^ m[796] ^ m[800] ^ m[805] ^ m[809] ^ m[810] ^ m[811] ^ m[815] ^ m[816] ^ m[817] ^ m[821] ^ m[822] ^ m[823] ^ m[827] ^ m[831] ^ m[832] ^ m[833] ^ m[837] ^ m[841] ^ m[846] ^ m[847] ^ m[848] ^ m[852] ^ m[856] ^ m[861] ^ m[867] ^ m[868] ^ m[869] ^ m[873] ^ m[877] ^ m[882] ^ m[888] ^ m[893] ^ m[894] ^ m[895] ^ m[899] ^ m[900] ^ m[901] ^ m[905] ^ m[906] ^ m[907] ^ m[911] ^ m[915] ^ m[916] ^ m[917] ^ m[921] ^ m[925] ^ m[930] ^ m[931] ^ m[932] ^ m[936] ^ m[940] ^ m[945] ^ m[951] ^ m[952] ^ m[953] ^ m[957] ^ m[961] ^ m[966] ^ m[972] ^ m[979] ^ m[980] ^ m[981] ^ m[985] ^ m[989] ^ m[994] ^ m[1000] ^ m[1007] ^ m[1012] ^ m[1013] ^ m[1014] ^ m[1015] ^ m[1017] ^ m[1018] ^ m[1019] ^ m[1020] ^ m[1021] ^ m[1022];
    assign parity[9] = m[0] ^ m[2] ^ m[3] ^ m[5] ^ m[6] ^ m[9] ^ m[11] ^ m[12] ^ m[15] ^ m[18] ^ m[21] ^ m[22] ^ m[25] ^ m[28] ^ m[32] ^ m[36] ^ m[37] ^ m[40] ^ m[43] ^ m[47] ^ m[52] ^ m[57] ^ m[58] ^ m[61] ^ m[64] ^ m[68] ^ m[73] ^ m[79] ^ m[85] ^ m[86] ^ m[89] ^ m[92] ^ m[96] ^ m[101] ^ m[107] ^ m[114] ^ m[121] ^ m[122] ^ m[125] ^ m[128] ^ m[132] ^ m[137] ^ m[143] ^ m[150] ^ m[158] ^ m[166] ^ m[167] ^ m[170] ^ m[173] ^ m[177] ^ m[182] ^ m[188] ^ m[195] ^ m[203] ^ m[212] ^ m[220] ^ m[221] ^ m[222] ^ m[224] ^ m[225] ^ m[226] ^ m[227] ^ m[229] ^ m[230] ^ m[231] ^ m[233] ^ m[234] ^ m[236] ^ m[237] ^ m[240] ^ m[241] ^ m[242] ^ m[244] ^ m[245] ^ m[246] ^ m[248] ^ m[249] ^ m[251] ^ m[252] ^ m[255] ^ m[256] ^ m[258] ^ m[259] ^ m[261] ^ m[262] ^ m[265] ^ m[267] ^ m[268] ^ m[271] ^ m[274] ^ m[276] ^ m[277] ^ m[279] ^ m[280] ^ m[281] ^ m[283] ^ m[284] ^ m[286] ^ m[287] ^ m[290] ^ m[291] ^ m[293] ^ m[294] ^ m[296] ^ m[297] ^ m[300] ^ m[302] ^ m[303] ^ m[306] ^ m[309] ^ m[311] ^ m[313] ^ m[314] ^ m[316] ^ m[317] ^ m[320] ^ m[322] ^ m[323] ^ m[326] ^ m[329] ^ m[332] ^ m[333] ^ m[336] ^ m[339] ^ m[343] ^ m[346] ^ m[347] ^ m[349] ^ m[350] ^ m[351] ^ m[353] ^ m[354] ^ m[356] ^ m[357] ^ m[360] ^ m[361] ^ m[363] ^ m[364] ^ m[366] ^ m[367] ^ m[370] ^ m[372] ^ m[373] ^ m[376] ^ m[379] ^ m[381] ^ m[383] ^ m[384] ^ m[386] ^ m[387] ^ m[390] ^ m[392] ^ m[393] ^ m[396] ^ m[399] ^ m[402] ^ m[403] ^ m[406] ^ m[409] ^ m[413] ^ m[416] ^ m[418] ^ m[419] ^ m[421] ^ m[422] ^ m[425] ^ m[427] ^ m[428] ^ m[431] ^ m[434] ^ m[437] ^ m[438] ^ m[441] ^ m[444] ^ m[448] ^ m[452] ^ m[453] ^ m[456] ^ m[459] ^ m[463] ^ m[468] ^ m[472] ^ m[473] ^ m[475] ^ m[476] ^ m[477] ^ m[479] ^ m[480] ^ m[482] ^ m[483] ^ m[486] ^ m[487] ^ m[489] ^ m[490] ^ m[492] ^ m[493] ^ m[496] ^ m[498] ^ m[499] ^ m[502] ^ m[505] ^ m[507] ^ m[509] ^ m[510] ^ m[512] ^ m[513] ^ m[516] ^ m[518] ^ m[519] ^ m[522] ^ m[525] ^ m[528] ^ m[529] ^ m[532] ^ m[535] ^ m[539] ^ m[542] ^ m[544] ^ m[545] ^ m[547] ^ m[548] ^ m[551] ^ m[553] ^ m[554] ^ m[557] ^ m[560] ^ m[563] ^ m[564] ^ m[567] ^ m[570] ^ m[574] ^ m[578] ^ m[579] ^ m[582] ^ m[585] ^ m[589] ^ m[594] ^ m[598] ^ m[600] ^ m[601] ^ m[603] ^ m[604] ^ m[607] ^ m[609] ^ m[610] ^ m[613] ^ m[616] ^ m[619] ^ m[620] ^ m[623] ^ m[626] ^ m[630] ^ m[634] ^ m[635] ^ m[638] ^ m[641] ^ m[645] ^ m[650] ^ m[655] ^ m[656] ^ m[659] ^ m[662] ^ m[666] ^ m[671] ^ m[677] ^ m[682] ^ m[683] ^ m[685] ^ m[686] ^ m[687] ^ m[689] ^ m[690] ^ m[692] ^ m[693] ^ m[696] ^ m[697] ^ m[699] ^ m[700] ^ m[702] ^ m[703] ^ m[706] ^ m[708] ^ m[709] ^ m[712] ^ m[715] ^ m[717] ^ m[719] ^ m[720] ^ m[722] ^ m[723] ^ m[726] ^ m[728] ^ m[729] ^ m[732] ^ m[735] ^ m[738] ^ m[739] ^ m[742] ^ m[745] ^ m[749] ^ m[752] ^ m[754] ^ m[755] ^ m[757] ^ m[758] ^ m[761] ^ m[763] ^ m[764] ^ m[767] ^ m[770] ^ m[773] ^ m[774] ^ m[777] ^ m[780] ^ m[784] ^ m[788] ^ m[789] ^ m[792] ^ m[795] ^ m[799] ^ m[804] ^ m[808] ^ m[810] ^ m[811] ^ m[813] ^ m[814] ^ m[817] ^ m[819] ^ m[820] ^ m[823] ^ m[826] ^ m[829] ^ m[830] ^ m[833] ^ m[836] ^ m[840] ^ m[844] ^ m[845] ^ m[848] ^ m[851] ^ m[855] ^ m[860] ^ m[865] ^ m[866] ^ m[869] ^ m[872] ^ m[876] ^ m[881] ^ m[887] ^ m[892] ^ m[894] ^ m[895] ^ m[897] ^ m[898] ^ m[901] ^ m[903] ^ m[904] ^ m[907] ^ m[910] ^ m[913] ^ m[914] ^ m[917] ^ m[920] ^ m[924] ^ m[928] ^ m[929] ^ m[932] ^ m[935] ^ m[939] ^ m[944] ^ m[949] ^ m[950] ^ m[953] ^ m[956] ^ m[960] ^ m[965] ^ m[971] ^ m[977] ^ m[978] ^ m[981] ^ m[984] ^ m[988] ^ m[993] ^ m[999] ^ m[1006] ^ m[1012] ^ m[1013] ^ m[1014] ^ m[1015] ^ m[1016] ^ m[1018] ^ m[1019] ^ m[1020] ^ m[1021] ^ m[1022] ^ m[1023];
    assign parity[10] = m[0] ^ m[1] ^ m[3] ^ m[4] ^ m[6] ^ m[8] ^ m[10] ^ m[12] ^ m[14] ^ m[17] ^ m[20] ^ m[22] ^ m[24] ^ m[27] ^ m[31] ^ m[35] ^ m[37] ^ m[39] ^ m[42] ^ m[46] ^ m[51] ^ m[56] ^ m[58] ^ m[60] ^ m[63] ^ m[67] ^ m[72] ^ m[78] ^ m[84] ^ m[86] ^ m[88] ^ m[91] ^ m[95] ^ m[100] ^ m[106] ^ m[113] ^ m[120] ^ m[122] ^ m[124] ^ m[127] ^ m[131] ^ m[136] ^ m[142] ^ m[149] ^ m[157] ^ m[165] ^ m[167] ^ m[169] ^ m[172] ^ m[176] ^ m[181] ^ m[187] ^ m[194] ^ m[202] ^ m[211] ^ m[220] ^ m[221] ^ m[222] ^ m[223] ^ m[225] ^ m[226] ^ m[227] ^ m[228] ^ m[230] ^ m[231] ^ m[232] ^ m[234] ^ m[235] ^ m[237] ^ m[239] ^ m[241] ^ m[242] ^ m[243] ^ m[245] ^ m[246] ^ m[247] ^ m[249] ^ m[250] ^ m[252] ^ m[254] ^ m[256] ^ m[257] ^ m[259] ^ m[260] ^ m[262] ^ m[264] ^ m[266] ^ m[268] ^ m[270] ^ m[273] ^ m[276] ^ m[277] ^ m[278] ^ m[280] ^ m[281] ^ m[282] ^ m[284] ^ m[285] ^ m[287] ^ m[289] ^ m[291] ^ m[292] ^ m[294] ^ m[295] ^ m[297] ^ m[299] ^ m[301] ^ m[303] ^ m[305] ^ m[308] ^ m[311] ^ m[312] ^ m[314] ^ m[315] ^ m[317] ^ m[319] ^ m[321] ^ m[323] ^ m[325] ^ m[328] ^ m[331] ^ m[333] ^ m[335] ^ m[338] ^ m[342] ^ m[346] ^ m[347] ^ m[348] ^ m[350] ^ m[351] ^ m[352] ^ m[354] ^ m[355] ^ m[357] ^ m[359] ^ m[361] ^ m[362] ^ m[364] ^ m[365] ^ m[367] ^ m[369] ^ m[371] ^ m[373] ^ m[375] ^ m[378] ^ m[381] ^ m[382] ^ m[384] ^ m[385] ^ m[387] ^ m[389] ^ m[391] ^ m[393] ^ m[395] ^ m[398] ^ m[401] ^ m[403] ^ m[405] ^ m[408] ^ m[412] ^ m[416] ^ m[417] ^ m[419] ^ m[420] ^ m[422] ^ m[424] ^ m[426] ^ m[428] ^ m[430] ^ m[433] ^ m[436] ^ m[438] ^ m[440] ^ m[443] ^ m[447] ^ m[451] ^ m[453] ^ m[455] ^ m[458] ^ m[462] ^ m[467] ^ m[472] ^ m[473] ^ m[474] ^ m[476] ^ m[477] ^ m[478] ^ m[480] ^ m[481] ^ m[483] ^ m[485] ^ m[487] ^ m[488] ^ m[490] ^ m[491] ^ m[493] ^ m[495] ^ m[497] ^ m[499] ^ m[501] ^ m[504] ^ m[507] ^ m[508] ^ m[510] ^ m[511] ^ m[513] ^ m[515] ^ m[517] ^ m[519] ^ m[521] ^ m[524] ^ m[527] ^ m[529] ^ m[531] ^ m[534] ^ m[538] ^ m[542] ^ m[543] ^ m[545] ^ m[546] ^ m[548] ^ m[550] ^ m[552] ^ m[554] ^ m[556] ^ m[559] ^ m[562] ^ m[564] ^ m[566] ^ m[569] ^ m[573] ^ m[577] ^ m[579] ^ m[581] ^ m[584] ^ m[588] ^ m[593] ^ m[598] ^ m[599] ^ m[601] ^ m[602] ^ m[604] ^ m[606] ^ m[608] ^ m[610] ^ m[612] ^ m[615] ^ m[618] ^ m[620] ^ m[622] ^ m[625] ^ m[629] ^ m[633] ^ m[635] ^ m[637] ^ m[640] ^ m[644] ^ m[649] ^ m[654] ^ m[656] ^ m[658] ^ m[661] ^ m[665] ^ m[670] ^ m[676] ^ m[682] ^ m[683] ^ m[684] ^ m[686] ^ m[687] ^ m[688] ^ m[690] ^ m[691] ^ m[693] ^ m[695] ^ m[697] ^ m[698] ^ m[700] ^ m[701] ^ m[703] ^ m[705] ^ m[707] ^ m[709] ^ m[711] ^ m[714] ^ m[717] ^ m[718] ^ m[720] ^ m[721] ^ m[723] ^ m[725] ^ m[727] ^ m[729] ^ m[731] ^ m[734] ^ m[737] ^ m[739] ^ m[741] ^ m[744] ^ m[748] ^ m[752] ^ m[753] ^ m[755] ^ m[756] ^ m[758] ^ m[760] ^ m[762] ^ m[764] ^ m[766] ^ m[769] ^ m[772] ^ m[774] ^ m[776] ^ m[779] ^ m[783] ^ m[787] ^ m[789] ^ m[791] ^ m[794] ^ m[798] ^ m[803] ^ m[808] ^ m[809] ^ m[811] ^ m[812] ^ m[814] ^ m[816] ^ m[818] ^ m[820] ^ m[822] ^ m[825] ^ m[828] ^ m[830] ^ m[832] ^ m[835] ^ m[839] ^ m[843] ^ m[845] ^ m[847] ^ m[850] ^ m[854] ^ m[859] ^ m[864] ^ m[866] ^ m[868] ^ m[871] ^ m[875] ^ m[880] ^ m[886] ^ m[892] ^ m[893] ^ m[895] ^ m[896] ^ m[898] ^ m[900] ^ m[902] ^ m[904] ^ m[906] ^ m[909] ^ m[912] ^ m[914] ^ m[916] ^ m[919] ^ m[923] ^ m[927] ^ m[929] ^ m[931] ^ m[934] ^ m[938] ^ m[943] ^ m[948] ^ m[950] ^ m[952] ^ m[955] ^ m[959] ^ m[964] ^ m[970] ^ m[976] ^ m[978] ^ m[980] ^ m[983] ^ m[987] ^ m[992] ^ m[998] ^ m[1005] ^ m[1012] ^ m[1013] ^ m[1014] ^ m[1015] ^ m[1016] ^ m[1017] ^ m[1019] ^ m[1020] ^ m[1021] ^ m[1022] ^ m[1023];
    assign parity[11] = m[0] ^ m[1] ^ m[2] ^ m[4] ^ m[5] ^ m[7] ^ m[10] ^ m[11] ^ m[13] ^ m[16] ^ m[20] ^ m[21] ^ m[23] ^ m[26] ^ m[30] ^ m[35] ^ m[36] ^ m[38] ^ m[41] ^ m[45] ^ m[50] ^ m[56] ^ m[57] ^ m[59] ^ m[62] ^ m[66] ^ m[71] ^ m[77] ^ m[84] ^ m[85] ^ m[87] ^ m[90] ^ m[94] ^ m[99] ^ m[105] ^ m[112] ^ m[120] ^ m[121] ^ m[123] ^ m[126] ^ m[130] ^ m[135] ^ m[141] ^ m[148] ^ m[156] ^ m[165] ^ m[166] ^ m[168] ^ m[171] ^ m[175] ^ m[180] ^ m[186] ^ m[193] ^ m[201] ^ m[210] ^ m[220] ^ m[221] ^ m[222] ^ m[223] ^ m[224] ^ m[226] ^ m[227] ^ m[228] ^ m[229] ^ m[231] ^ m[232] ^ m[233] ^ m[235] ^ m[236] ^ m[238] ^ m[241] ^ m[242] ^ m[243] ^ m[244] ^ m[246] ^ m[247] ^ m[248] ^ m[250] ^ m[251] ^ m[253] ^ m[256] ^ m[257] ^ m[258] ^ m[260] ^ m[261] ^ m[263] ^ m[266] ^ m[267] ^ m[269] ^ m[272] ^ m[276] ^ m[277] ^ m[278] ^ m[279] ^ m[281] ^ m[282] ^ m[283] ^ m[285] ^ m[286] ^ m[288] ^ m[291] ^ m[292] ^ m[293] ^ m[295] ^ m[296] ^ m[298] ^ m[301] ^ m[302] ^ m[304] ^ m[307] ^ m[311] ^ m[312] ^ m[313] ^ m[315] ^ m[316] ^ m[318] ^ m[321] ^ m[322] ^ m[324] ^ m[327] ^ m[331] ^ m[332] ^ m[334] ^ m[337] ^ m[341] ^ m[346] ^ m[347] ^ m[348] ^ m[349] ^ m[351] ^ m[352] ^ m[353] ^ m[355] ^ m[356] ^ m[358] ^ m[361] ^ m[362] ^ m[363] ^ m[365] ^ m[366] ^ m[368] ^ m[371] ^ m[372] ^ m[374] ^ m[377] ^ m[381] ^ m[382] ^ m[383] ^ m[385] ^ m[386] ^ m[388] ^ m[391] ^ m[392] ^ m[394] ^ m[397] ^ m[401] ^ m[402] ^ m[404] ^ m[407] ^ m[411] ^ m[416] ^ m[417] ^ m[418] ^ m[420] ^ m[421] ^ m[423] ^ m[426] ^ m[427] ^ m[429] ^ m[432] ^ m[436] ^ m[437] ^ m[439] ^ m[442] ^ m[446] ^ m[451] ^ m[452] ^ m[454] ^ m[457] ^ m[461] ^ m[466] ^ m[472] ^ m[473] ^ m[474] ^ m[475] ^ m[477] ^ m[478] ^ m[479] ^ m[481] ^ m[482] ^ m[484] ^ m[487] ^ m[488] ^ m[489] ^ m[491] ^ m[492] ^ m[494] ^ m[497] ^ m[498] ^ m[500] ^ m[503] ^ m[507] ^ m[508] ^ m[509] ^ m[511] ^ m[512] ^ m[514] ^ m[517] ^ m[518] ^ m[520] ^ m[523] ^ m[527] ^ m[528] ^ m[530] ^ m[533] ^ m[537] ^ m[542] ^ m[543] ^ m[544] ^ m[546] ^ m[547] ^ m[549] ^ m[552] ^ m[553] ^ m[555] ^ m[558] ^ m[562] ^ m[563] ^ m[565] ^ m[568] ^ m[572] ^ m[577] ^ m[578] ^ m[580] ^ m[583] ^ m[587] ^ m[592] ^ m[598] ^ m[599] ^ m[600] ^ m[602] ^ m[603] ^ m[605] ^ m[608] ^ m[609] ^ m[611] ^ m[614] ^ m[618] ^ m[619] ^ m[621] ^ m[624] ^ m[628] ^ m[633] ^ m[634] ^ m[636] ^ m[639] ^ m[643] ^ m[648] ^ m[654] ^ m[655] ^ m[657] ^ m[660] ^ m[664] ^ m[669] ^ m[675] ^ m[682] ^ m[683] ^ m[684] ^ m[685] ^ m[687] ^ m[688] ^ m[689] ^ m[691] ^ m[692] ^ m[694] ^ m[697] ^ m[698] ^ m[699] ^ m[701] ^ m[702] ^ m[704] ^ m[707] ^ m[708] ^ m[710] ^ m[713] ^ m[717] ^ m[718] ^ m[719] ^ m[721] ^ m[722] ^ m[724] ^ m[727] ^ m[728] ^ m[730] ^ m[733] ^ m[737] ^ m[738] ^ m[740] ^ m[743] ^ m[747] ^ m[752] ^ m[753] ^ m[754] ^ m[756] ^ m[757] ^ m[759] ^ m[762] ^ m[763] ^ m[765] ^ m[768] ^ m[772] ^ m[773] ^ m[775] ^ m[778] ^ m[782] ^ m[787] ^ m[788] ^ m[790] ^ m[793] ^ m[797] ^ m[802] ^ m[808] ^ m[809] ^ m[810] ^ m[812] ^ m[813] ^ m[815] ^ m[818] ^ m[819] ^ m[821] ^ m[824] ^ m[828] ^ m[829] ^ m[831] ^ m[834] ^ m[838] ^ m[843] ^ m[844] ^ m[846] ^ m[849] ^ m[853] ^ m[858] ^ m[864] ^ m[865] ^ m[867] ^ m[870] ^ m[874] ^ m[879] ^ m[885] ^ m[892] ^ m[893] ^ m[894] ^ m[896] ^ m[897] ^ m[899] ^ m[902] ^ m[903] ^ m[905] ^ m[908] ^ m[912] ^ m[913] ^ m[915] ^ m[918] ^ m[922] ^ m[927] ^ m[928] ^ m[930] ^ m[933] ^ m[937] ^ m[942] ^ m[948] ^ m[949] ^ m[951] ^ m[954] ^ m[958] ^ m[963] ^ m[969] ^ m[976] ^ m[977] ^ m[979] ^ m[982] ^ m[986] ^ m[991] ^ m[997] ^ m[1004] ^ m[1012] ^ m[1013] ^ m[1014] ^ m[1015] ^ m[1016] ^ m[1017] ^ m[1018] ^ m[1020] ^ m[1021] ^ m[1022] ^ m[1023];
  end else begin : gen_default_parity
    `BR_ASSERT_STATIC(invalid_parity_width_a, 1'b0)
  end

  // ri lint_check_on EXPR_ID_LIMIT

  //------
  // Concatenate message and parity bits to form the codeword.
  //------
  logic [CodewordWidth-1:0] internal_codeword;
  assign internal_codeword = {parity, m};

  //------
  // Optionally register the output signals.
  //------
  br_delay_valid #(
      .Width(CodewordWidth),
      .NumStages(RegisterOutputs == 1 ? 1 : 0)
  ) br_delay_valid_outputs (
      .clk,
      .rst,
      .in_valid(data_valid_d),
      .in({internal_codeword}),
      .out_valid(enc_valid),
      .out(enc_codeword),
      .out_valid_stages(),  // unused
      .out_stages()  // unused
  );

  //------------------------------------------
  // Implementation checks
  //------------------------------------------
  `BR_ASSERT_IMPL(latency_a, data_valid |-> ##Latency enc_valid)

  // verilog_lint: waive-stop line-length
  // verilog_format: on

endmodule : br_ecc_secded_encoder
