// Copyright 2024 The Bedrock-RTL Authors
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//     http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.

`include "br_asserts_internal.svh"
`include "br_registers.svh"

module br_credit_sender #(
    // Width of the datapath in bits. Must be at least 1.
    parameter int BitWidth = 1,
    // Maximum number of credits that can be stored (inclusive). Must be at least 1.
    parameter int MaxCredit = 1,
    localparam int CounterWidth = $clog2(MaxCredit + 1)
) (
    // Posedge-triggered clock.
    input logic clk,
    // Synchronous active-high reset.
    input logic rst,
    input logic [CounterWidth-1:0] initial_credit,
    // Ready/valid push interface.
    output logic push_ready,
    input logic push_valid,
    input logic [BitWidth-1:0] push_data,
    // Credit/valid pop interface.
    output logic pop_credit_stall,
    input logic pop_credit,
    output logic pop_valid,
    output logic [BitWidth-1:0] pop_data,
    output logic [CounterWidth-1:0] credit_count
);

  //------------------------------------------
  // Integration checks
  //------------------------------------------
  `BR_ASSERT_STATIC(bitwidth_in_range_a, BitWidth >= 1)
  `BR_ASSERT_STATIC(max_credit_in_range_a, MaxCredit >= 1)

  `BR_ASSERT_INTG(no_pop_credit_when_stall_a, pop_credit_stall |-> !pop_credit)

  // TODO(mgottscho): write some

  //------------------------------------------
  // Implementation
  //------------------------------------------
  br_credit_counter #(
      .MaxValue (MaxCredit),
      .MaxChange(1)
  ) br_credit_counter (
      .clk,
      .rst,
      .initial_value(initial_credit),
      .incr_valid(pop_credit),
      .incr(1'b1),
      .decr_valid(pop_valid),
      .decr(1'b1),
      .value(credit_count),
      .value_next()  // unused
  );

  `BR_REGI(pop_credit_stall, 1'b0, 1'b1);
  assign push_ready = credit_count > 0;
  assign pop_valid  = push_ready && push_valid;
  assign pop_data   = push_data;

  //------------------------------------------
  // Implementation checks
  //------------------------------------------

  // TODO(mgottscho): write some

endmodule : br_credit_sender
