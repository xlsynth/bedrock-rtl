// Copyright 2024 The Bedrock-RTL Authors
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//     http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.

// Bedrock-RTL Incrementing Counter
//
// A simple counter that increments by a potentially variable amount each cycle,
// where the maximum increment is given by MaxIncrement (inclusive).
// Overflows (wraps around past 0) at MaxValue (inclusive), even if MaxValue + 1
// isn't a power-of-2. In the common case where MaxValue + 1 is a power-of-2,
// the implementation is simplified.
//
// When there is a valid increment and it overflows:
//   value_next = (value + incr) % (MaxValue + 1)
//
// The counter state is exposed in two ways.
// (1) value holds the current counter state. There is a latency of 1 cycle from
//     a valid increment to the counter state being updated.
// (2) value_next is what value will be on the next cycle. It is conditioned on
//     incr_valid: if low, then value_next == value. This is useful for constructing
//     single-cycle chains of counters.
// value and value_next are always valid.
//
// The value resets to 0.

`include "br_asserts_internal.svh"
`include "br_registers.svh"

module br_counter_incr #(
    parameter int MaxValue = 1,  // Must be at least 1. Inclusive.
    parameter int MaxIncrement = 1,  // Must be at least 1 and at most MaxValue. Inclusive.
    localparam int ValueWidth = $clog2(MaxValue + 1),
    localparam int IncrementWidth = $clog2(MaxIncrement + 1)
) (
    input  logic                      clk,
    input  logic                      rst,
    input  logic                      incr_valid,
    input  logic [IncrementWidth-1:0] incr,
    output logic [    ValueWidth-1:0] value,
    output logic [    ValueWidth-1:0] value_next
);

  //------------------------------------------
  // Integration checks
  //------------------------------------------
  `BR_ASSERT_STATIC(max_value_gte_1_a, MaxValue >= 1)
  `BR_ASSERT_STATIC(max_increment_gte_1_a, MaxIncrement >= 1)
  `BR_ASSERT_STATIC(max_increment_lte_max_value_a, MaxIncrement <= MaxValue)

  `BR_ASSERT_INTG(incr_in_range_a, incr_valid |-> incr <= MaxIncrement)

  //------------------------------------------
  // Implementation
  //------------------------------------------
  localparam int MaxValueP1 = MaxValue + 1;
  localparam bit IsMaxValueP1PowerOf2 = (MaxValueP1 & (MaxValueP1 - 1)) == 0;
  localparam int TempWidth = $clog2(MaxValue + MaxIncrement + 1);

  logic [ValueWidth-1:0] value_next_internal;

  // TODO(mgottscho): Sometimes the MSbs may not be used. It'd be cleaner
  // to capture them more tightly using br_misc_unused.
  // ri lint_check_waive NOT_READ
  logic [ TempWidth-1:0] value_temp;
  assign value_temp = value + incr;

  // For MaxValueP1 being a power of 2, wrapping occurs naturally
  if (IsMaxValueP1PowerOf2) begin : gen_power_of_2
    assign value_next_internal = incr_valid ? value_temp[ValueWidth-1:0] : value;

    // For MaxValueP1 not being a power of 2, handle wrap-around explicitly
  end else begin : gen_non_power_of_2
    // MSBs won't impact outputs if TempWidth > ValueWidth
    // ri lint_check_waive INEFFECTIVE_NET
    logic [TempWidth-1:0] value_temp_wrapped;

    // ri lint_check_waive ARITH_EXTENSION
    assign value_temp_wrapped = (value_temp - MaxValue) - 1;
    // ri lint_check_waive ARITH_EXTENSION
    assign value_next_internal = (value_temp >= MaxValue) ?
      value_temp_wrapped[ValueWidth-1:0] :  // ri lint_check_waive FULL_RANGE
        value_temp[ValueWidth-1:0];  // ri lint_check_waive FULL_RANGE

    if (TempWidth > ValueWidth) begin : gen_unused
      br_misc_unused #(
          .BitWidth(TempWidth - ValueWidth)
      ) br_misc_unused_value_temp_wrapped_msbs (
          .in(value_temp_wrapped[TempWidth-1:ValueWidth])
      );
    end
  end

  // If the user leaves the value_next port unused, then the synthesis tool
  // should be able to automatically simplify the following ternary expression
  // to just value_next_internal, because the load-enable on the register is
  // conditioned on the same incr_valid.
  assign value_next = incr_valid ? value_next_internal : value;
  `BR_REGL(value, value_next, incr_valid)

  //------------------------------------------
  // Implementation checks
  //------------------------------------------
  `BR_ASSERT_IMPL(value_in_range_a, value <= MaxValue)
  `BR_ASSERT_IMPL(value_next_in_range_a, value_next <= MaxValue)
  `BR_ASSERT_IMPL(value_next_propagates_a, ##1 value == $past(value_next))
  `BR_ASSERT_IMPL(value_wrap_a,
                  incr_valid && value_temp > MaxValue |-> value_next == value_temp - MaxValue - 1)
  `BR_ASSERT_IMPL(maxvalue_plus_one_a,
                  value == MaxValue && incr_valid && incr == 1'b1 |-> value_next == 0)
  `BR_ASSERT_IMPL(plus_zero_a, incr_valid && incr == '0 |-> value_next == value)
  `BR_COVER_IMPL(increment_max_c, incr_valid && incr == MaxIncrement)
  `BR_COVER_IMPL(value_temp_oob_c, value_temp > MaxValue)

endmodule : br_counter_incr
