// Copyright 2024 The Bedrock-RTL Authors
//
// Licensed under the Apache License, Version 2.0 (the "License");
// Copyright 2024 The Bedrock-RTL Authors
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//     http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.


// verilog_format: off
// verilog_lint: waive-start line-length

// Bedrock-RTL Single-Error-Correcting, Double-Error-Detecting (SECDED - Hsiao) Encoder
//
// Encodes a message using a single-error-correcting, double-error-detecting
// linear block code in systematic form (in layperson's terms: a Hsiao SECDED [1] encoder,
// closely related to Hamming codes).
//
// Systematic form means that the codeword is formed by appending the
// calculated parity bits to the message, i.e., the code has the property
// that the message bits are 1:1 with a slice of bits in the codeword (if they
// have not been corrupted).
//
// In Bedrock ECC libs, our convention is to always append the parity bits on
// the MSbs:
//     codeword == {parity, message}
//
// This module has a parameterizable number of pipeline stages, ranging from fully
// combinational to 1 cycle of latency.
//
// Any data width >= 1 is supported. It is internally zero-padded up to
// the nearest power-of-2 message width before being encoded. The following
// table outlines the number of parity bits required for different message widths.
//
// | Message Width (k) | Parity Width (r) | Codeword Width (n)|
// |-------------------|------------------|-------------------|
// | 4                 | 4                | 8                 |
// | 8                 | 5                | 13                |
// | 16                | 6                | 22                |
// | 32                | 7                | 39                |
// | 64                | 8                | 72                |
// | 128               | 9                | 137               |
// | 256               | 10               | 266               |
// | 512               | 11               | 523               |
// | 1024              | 12               | 1036              |
//
// The number of parity bits must be one of the values in the table above
// or the module will not elaborate.
//
// References:
// [1] https://ieeexplore.ieee.org/abstract/document/5391627

`include "br_asserts.svh"
`include "br_asserts_internal.svh"

module br_ecc_secded_encoder #(
    parameter int DataWidth = 1,  // Must be at least 1
    parameter int ParityWidth = 4,  // Must be at least 4 and at most 12
    // If 1, then insert a pipeline register at the output.
    parameter bit RegisterOutputs = 0,
    localparam int MessageWidth = 2 ** $clog2(DataWidth),
    localparam int CodewordWidth = MessageWidth + ParityWidth
) (
    // Positive edge-triggered clock.
    input  logic                     clk,
    // Synchronous active-high reset.
    input  logic                     rst,
    input  logic                     data_valid,
    input  logic [    DataWidth-1:0] data,
    output logic                     codeword_valid,
    output logic [CodewordWidth-1:0] codeword
);

  // ri lint_check_waive PARAM_NOT_USED
  localparam int Latency = RegisterOutputs ? 1 : 0;

  //------------------------------------------
  // Integration checks
  //------------------------------------------
  `BR_ASSERT_STATIC(message_width_gte_1_a, DataWidth >= 1)
  `BR_ASSERT_STATIC(parity_width_gte_4_a, ParityWidth >= 4)
  `BR_ASSERT_STATIC(parity_width_lte_12_a, ParityWidth <= 12)
  `BR_ASSERT_STATIC(message_width_is_power_of_2_a, br_math::is_power_of_2(MessageWidth))

  //------------------------------------------
  // Implementation
  //------------------------------------------


  //------
  // Pad data to the nearest power of 2 message width.
  //------
  localparam int PadWidth = MessageWidth - DataWidth;
  logic [MessageWidth-1:0] message;

  if (PadWidth > 0) begin : gen_pad
    assign message = { {PadWidth{1'b0} }, data};
  end else begin : gen_no_pad
    assign message = data;
  end

  //------
  // Compute parity bits.
  //------
  logic [ParityWidth-1:0] parity;

  // ri lint_check_off EXPR_ID_LIMIT

  if ((CodewordWidth == 4) && (MessageWidth == 4)) begin : gen_8_4
    `BR_ASSERT_STATIC(parity_width_matches_a, ParityWidth == 4)
    assign parity[0] = message[1] ^ message[2] ^ message[3];
    assign parity[1] = message[0] ^ message[2] ^ message[3];
    assign parity[2] = message[0] ^ message[1] ^ message[3];
    assign parity[3] = message[0] ^ message[1] ^ message[2];
  end else if ((CodewordWidth == 13) && (MessageWidth == 8)) begin : gen_13_8
    `BR_ASSERT_STATIC(parity_width_matches_a, ParityWidth == 5)
    assign parity[0] = message[4] ^ message[5] ^ message[6] ^ message[7];
    assign parity[1] = message[1] ^ message[2] ^ message[3] ^ message[7];
    assign parity[2] = message[0] ^ message[2] ^ message[3] ^ message[5] ^ message[6];
    assign parity[3] = message[0] ^ message[1] ^ message[3] ^ message[4] ^ message[6];
    assign parity[4] = message[0] ^ message[1] ^ message[2] ^ message[4] ^ message[5] ^ message[7];
  end else if ((CodewordWidth == 22) && (MessageWidth == 16)) begin : gen_22_16
    `BR_ASSERT_STATIC(parity_width_matches_a, ParityWidth == 6)
    assign parity[0] = message[10] ^ message[11] ^ message[12] ^ message[13] ^ message[14] ^ message[15];
    assign parity[1] = message[4] ^ message[5] ^ message[6] ^ message[7] ^ message[8] ^ message[9];
    assign parity[2] = message[1] ^ message[2] ^ message[3] ^ message[7] ^ message[8] ^ message[9] ^ message[13] ^ message[14] ^ message[15];
    assign parity[3] = message[0] ^ message[2] ^ message[3] ^ message[5] ^ message[6] ^ message[9] ^ message[11] ^ message[12] ^ message[15];
    assign parity[4] = message[0] ^ message[1] ^ message[3] ^ message[4] ^ message[6] ^ message[8] ^ message[10] ^ message[12] ^ message[14];
    assign parity[5] = message[0] ^ message[1] ^ message[2] ^ message[4] ^ message[5] ^ message[7] ^ message[10] ^ message[11] ^ message[13];
  end else if ((CodewordWidth == 39) && (MessageWidth == 32)) begin : gen_39_32
    `BR_ASSERT_STATIC(parity_width_matches_a, ParityWidth == 7)
    assign parity[0] = message[20] ^ message[21] ^ message[22] ^ message[23] ^ message[24] ^ message[25] ^ message[26] ^ message[27] ^ message[28] ^ message[29] ^ message[30] ^ message[31];
    assign parity[1] = message[10] ^ message[11] ^ message[12] ^ message[13] ^ message[14] ^ message[15] ^ message[16] ^ message[17] ^ message[18] ^ message[19] ^ message[30] ^ message[31];
    assign parity[2] = message[4] ^ message[5] ^ message[6] ^ message[7] ^ message[8] ^ message[9] ^ message[16] ^ message[17] ^ message[18] ^ message[19] ^ message[26] ^ message[27] ^ message[28] ^ message[29];
    assign parity[3] = message[1] ^ message[2] ^ message[3] ^ message[7] ^ message[8] ^ message[9] ^ message[13] ^ message[14] ^ message[15] ^ message[19] ^ message[23] ^ message[24] ^ message[25] ^ message[29];
    assign parity[4] = message[0] ^ message[2] ^ message[3] ^ message[5] ^ message[6] ^ message[9] ^ message[11] ^ message[12] ^ message[15] ^ message[18] ^ message[21] ^ message[22] ^ message[25] ^ message[28];
    assign parity[5] = message[0] ^ message[1] ^ message[3] ^ message[4] ^ message[6] ^ message[8] ^ message[10] ^ message[12] ^ message[14] ^ message[17] ^ message[20] ^ message[22] ^ message[24] ^ message[27] ^ message[31];
    assign parity[6] = message[0] ^ message[1] ^ message[2] ^ message[4] ^ message[5] ^ message[7] ^ message[10] ^ message[11] ^ message[13] ^ message[16] ^ message[20] ^ message[21] ^ message[23] ^ message[26] ^ message[30];
  end else if ((CodewordWidth == 72) && (MessageWidth == 64)) begin : gen_72_64
    `BR_ASSERT_STATIC(parity_width_matches_a, ParityWidth == 8)
    assign parity[0] = message[35] ^ message[36] ^ message[37] ^ message[38] ^ message[39] ^ message[40] ^ message[41] ^ message[42] ^ message[43] ^ message[44] ^ message[45] ^ message[46] ^ message[47] ^ message[48] ^ message[49] ^ message[50] ^ message[51] ^ message[52] ^ message[53] ^ message[54] ^ message[55];
    assign parity[1] = message[20] ^ message[21] ^ message[22] ^ message[23] ^ message[24] ^ message[25] ^ message[26] ^ message[27] ^ message[28] ^ message[29] ^ message[30] ^ message[31] ^ message[32] ^ message[33] ^ message[34] ^ message[50] ^ message[51] ^ message[52] ^ message[53] ^ message[54] ^ message[55] ^ message[62] ^ message[63];
    assign parity[2] = message[10] ^ message[11] ^ message[12] ^ message[13] ^ message[14] ^ message[15] ^ message[16] ^ message[17] ^ message[18] ^ message[19] ^ message[30] ^ message[31] ^ message[32] ^ message[33] ^ message[34] ^ message[45] ^ message[46] ^ message[47] ^ message[48] ^ message[49] ^ message[55] ^ message[57] ^ message[58] ^ message[59] ^ message[60] ^ message[61];
    assign parity[3] = message[4] ^ message[5] ^ message[6] ^ message[7] ^ message[8] ^ message[9] ^ message[16] ^ message[17] ^ message[18] ^ message[19] ^ message[26] ^ message[27] ^ message[28] ^ message[29] ^ message[34] ^ message[41] ^ message[42] ^ message[43] ^ message[44] ^ message[49] ^ message[54] ^ message[56] ^ message[58] ^ message[59] ^ message[60] ^ message[61] ^ message[63];
    assign parity[4] = message[1] ^ message[2] ^ message[3] ^ message[7] ^ message[8] ^ message[9] ^ message[13] ^ message[14] ^ message[15] ^ message[19] ^ message[23] ^ message[24] ^ message[25] ^ message[29] ^ message[33] ^ message[38] ^ message[39] ^ message[40] ^ message[44] ^ message[48] ^ message[53] ^ message[56] ^ message[57] ^ message[59] ^ message[60] ^ message[61] ^ message[62];
    assign parity[5] = message[0] ^ message[2] ^ message[3] ^ message[5] ^ message[6] ^ message[9] ^ message[11] ^ message[12] ^ message[15] ^ message[18] ^ message[21] ^ message[22] ^ message[25] ^ message[28] ^ message[32] ^ message[36] ^ message[37] ^ message[40] ^ message[43] ^ message[47] ^ message[52] ^ message[56] ^ message[57] ^ message[58] ^ message[60] ^ message[61] ^ message[62] ^ message[63];
    assign parity[6] = message[0] ^ message[1] ^ message[3] ^ message[4] ^ message[6] ^ message[8] ^ message[10] ^ message[12] ^ message[14] ^ message[17] ^ message[20] ^ message[22] ^ message[24] ^ message[27] ^ message[31] ^ message[35] ^ message[37] ^ message[39] ^ message[42] ^ message[46] ^ message[51] ^ message[56] ^ message[57] ^ message[58] ^ message[59] ^ message[61] ^ message[62] ^ message[63];
    assign parity[7] = message[0] ^ message[1] ^ message[2] ^ message[4] ^ message[5] ^ message[7] ^ message[10] ^ message[11] ^ message[13] ^ message[16] ^ message[20] ^ message[21] ^ message[23] ^ message[26] ^ message[30] ^ message[35] ^ message[36] ^ message[38] ^ message[41] ^ message[45] ^ message[50] ^ message[56] ^ message[57] ^ message[58] ^ message[59] ^ message[60] ^ message[62] ^ message[63];
  end else if ((CodewordWidth == 137) && (MessageWidth == 128)) begin : gen_137_128
    `BR_ASSERT_STATIC(parity_width_matches_a, ParityWidth == 9)
    assign parity[0] = message[56] ^ message[57] ^ message[58] ^ message[59] ^ message[60] ^ message[61] ^ message[62] ^ message[63] ^ message[64] ^ message[65] ^ message[66] ^ message[67] ^ message[68] ^ message[69] ^ message[70] ^ message[71] ^ message[72] ^ message[73] ^ message[74] ^ message[75] ^ message[76] ^ message[77] ^ message[78] ^ message[79] ^ message[80] ^ message[81] ^ message[82] ^ message[83];
    assign parity[1] = message[35] ^ message[36] ^ message[37] ^ message[38] ^ message[39] ^ message[40] ^ message[41] ^ message[42] ^ message[43] ^ message[44] ^ message[45] ^ message[46] ^ message[47] ^ message[48] ^ message[49] ^ message[50] ^ message[51] ^ message[52] ^ message[53] ^ message[54] ^ message[55] ^ message[77] ^ message[78] ^ message[79] ^ message[80] ^ message[81] ^ message[82] ^ message[83] ^ message[105] ^ message[106] ^ message[107] ^ message[108] ^ message[109] ^ message[110] ^ message[111] ^ message[112] ^ message[113] ^ message[114] ^ message[115] ^ message[116] ^ message[117] ^ message[118] ^ message[119] ^ message[120] ^ message[121] ^ message[122] ^ message[123] ^ message[124] ^ message[125] ^ message[126] ^ message[127];
    assign parity[2] = message[20] ^ message[21] ^ message[22] ^ message[23] ^ message[24] ^ message[25] ^ message[26] ^ message[27] ^ message[28] ^ message[29] ^ message[30] ^ message[31] ^ message[32] ^ message[33] ^ message[34] ^ message[50] ^ message[51] ^ message[52] ^ message[53] ^ message[54] ^ message[55] ^ message[71] ^ message[72] ^ message[73] ^ message[74] ^ message[75] ^ message[76] ^ message[83] ^ message[90] ^ message[91] ^ message[92] ^ message[93] ^ message[94] ^ message[95] ^ message[96] ^ message[97] ^ message[98] ^ message[99] ^ message[100] ^ message[101] ^ message[102] ^ message[103] ^ message[104] ^ message[120] ^ message[121] ^ message[122] ^ message[123] ^ message[124] ^ message[125] ^ message[126] ^ message[127];
    assign parity[3] = message[10] ^ message[11] ^ message[12] ^ message[13] ^ message[14] ^ message[15] ^ message[16] ^ message[17] ^ message[18] ^ message[19] ^ message[30] ^ message[31] ^ message[32] ^ message[33] ^ message[34] ^ message[45] ^ message[46] ^ message[47] ^ message[48] ^ message[49] ^ message[55] ^ message[66] ^ message[67] ^ message[68] ^ message[69] ^ message[70] ^ message[76] ^ message[82] ^ message[85] ^ message[86] ^ message[87] ^ message[88] ^ message[89] ^ message[95] ^ message[96] ^ message[97] ^ message[98] ^ message[99] ^ message[100] ^ message[101] ^ message[102] ^ message[103] ^ message[104] ^ message[110] ^ message[111] ^ message[112] ^ message[113] ^ message[114] ^ message[115] ^ message[116] ^ message[117] ^ message[118] ^ message[119];
    assign parity[4] = message[4] ^ message[5] ^ message[6] ^ message[7] ^ message[8] ^ message[9] ^ message[16] ^ message[17] ^ message[18] ^ message[19] ^ message[26] ^ message[27] ^ message[28] ^ message[29] ^ message[34] ^ message[41] ^ message[42] ^ message[43] ^ message[44] ^ message[49] ^ message[54] ^ message[62] ^ message[63] ^ message[64] ^ message[65] ^ message[70] ^ message[75] ^ message[81] ^ message[84] ^ message[86] ^ message[87] ^ message[88] ^ message[89] ^ message[91] ^ message[92] ^ message[93] ^ message[94] ^ message[99] ^ message[100] ^ message[101] ^ message[102] ^ message[103] ^ message[104] ^ message[106] ^ message[107] ^ message[108] ^ message[109] ^ message[114] ^ message[115] ^ message[116] ^ message[117] ^ message[118] ^ message[119] ^ message[124] ^ message[125] ^ message[126] ^ message[127];
    assign parity[5] = message[1] ^ message[2] ^ message[3] ^ message[7] ^ message[8] ^ message[9] ^ message[13] ^ message[14] ^ message[15] ^ message[19] ^ message[23] ^ message[24] ^ message[25] ^ message[29] ^ message[33] ^ message[38] ^ message[39] ^ message[40] ^ message[44] ^ message[48] ^ message[53] ^ message[59] ^ message[60] ^ message[61] ^ message[65] ^ message[69] ^ message[74] ^ message[80] ^ message[84] ^ message[85] ^ message[87] ^ message[88] ^ message[89] ^ message[90] ^ message[92] ^ message[93] ^ message[94] ^ message[96] ^ message[97] ^ message[98] ^ message[102] ^ message[103] ^ message[104] ^ message[105] ^ message[107] ^ message[108] ^ message[109] ^ message[111] ^ message[112] ^ message[113] ^ message[117] ^ message[118] ^ message[119] ^ message[121] ^ message[122] ^ message[123] ^ message[127];
    assign parity[6] = message[0] ^ message[2] ^ message[3] ^ message[5] ^ message[6] ^ message[9] ^ message[11] ^ message[12] ^ message[15] ^ message[18] ^ message[21] ^ message[22] ^ message[25] ^ message[28] ^ message[32] ^ message[36] ^ message[37] ^ message[40] ^ message[43] ^ message[47] ^ message[52] ^ message[57] ^ message[58] ^ message[61] ^ message[64] ^ message[68] ^ message[73] ^ message[79] ^ message[84] ^ message[85] ^ message[86] ^ message[88] ^ message[89] ^ message[90] ^ message[91] ^ message[93] ^ message[94] ^ message[95] ^ message[97] ^ message[98] ^ message[100] ^ message[101] ^ message[104] ^ message[105] ^ message[106] ^ message[108] ^ message[109] ^ message[110] ^ message[112] ^ message[113] ^ message[115] ^ message[116] ^ message[119] ^ message[120] ^ message[122] ^ message[123] ^ message[125] ^ message[126];
    assign parity[7] = message[0] ^ message[1] ^ message[3] ^ message[4] ^ message[6] ^ message[8] ^ message[10] ^ message[12] ^ message[14] ^ message[17] ^ message[20] ^ message[22] ^ message[24] ^ message[27] ^ message[31] ^ message[35] ^ message[37] ^ message[39] ^ message[42] ^ message[46] ^ message[51] ^ message[56] ^ message[58] ^ message[60] ^ message[63] ^ message[67] ^ message[72] ^ message[78] ^ message[84] ^ message[85] ^ message[86] ^ message[87] ^ message[89] ^ message[90] ^ message[91] ^ message[92] ^ message[94] ^ message[95] ^ message[96] ^ message[98] ^ message[99] ^ message[101] ^ message[103] ^ message[105] ^ message[106] ^ message[107] ^ message[109] ^ message[110] ^ message[111] ^ message[113] ^ message[114] ^ message[116] ^ message[118] ^ message[120] ^ message[121] ^ message[123] ^ message[124] ^ message[126];
    assign parity[8] = message[0] ^ message[1] ^ message[2] ^ message[4] ^ message[5] ^ message[7] ^ message[10] ^ message[11] ^ message[13] ^ message[16] ^ message[20] ^ message[21] ^ message[23] ^ message[26] ^ message[30] ^ message[35] ^ message[36] ^ message[38] ^ message[41] ^ message[45] ^ message[50] ^ message[56] ^ message[57] ^ message[59] ^ message[62] ^ message[66] ^ message[71] ^ message[77] ^ message[84] ^ message[85] ^ message[86] ^ message[87] ^ message[88] ^ message[90] ^ message[91] ^ message[92] ^ message[93] ^ message[95] ^ message[96] ^ message[97] ^ message[99] ^ message[100] ^ message[102] ^ message[105] ^ message[106] ^ message[107] ^ message[108] ^ message[110] ^ message[111] ^ message[112] ^ message[114] ^ message[115] ^ message[117] ^ message[120] ^ message[121] ^ message[122] ^ message[124] ^ message[125] ^ message[127];
  end else if ((CodewordWidth == 266) && (MessageWidth == 256)) begin : gen_266_256
    `BR_ASSERT_STATIC(parity_width_matches_a, ParityWidth == 10)
    assign parity[0] = message[84] ^ message[85] ^ message[86] ^ message[87] ^ message[88] ^ message[89] ^ message[90] ^ message[91] ^ message[92] ^ message[93] ^ message[94] ^ message[95] ^ message[96] ^ message[97] ^ message[98] ^ message[99] ^ message[100] ^ message[101] ^ message[102] ^ message[103] ^ message[104] ^ message[105] ^ message[106] ^ message[107] ^ message[108] ^ message[109] ^ message[110] ^ message[111] ^ message[112] ^ message[113] ^ message[114] ^ message[115] ^ message[116] ^ message[117] ^ message[118] ^ message[119] ^ message[246] ^ message[247] ^ message[248] ^ message[249] ^ message[250] ^ message[251] ^ message[252] ^ message[253] ^ message[254] ^ message[255];
    assign parity[1] = message[56] ^ message[57] ^ message[58] ^ message[59] ^ message[60] ^ message[61] ^ message[62] ^ message[63] ^ message[64] ^ message[65] ^ message[66] ^ message[67] ^ message[68] ^ message[69] ^ message[70] ^ message[71] ^ message[72] ^ message[73] ^ message[74] ^ message[75] ^ message[76] ^ message[77] ^ message[78] ^ message[79] ^ message[80] ^ message[81] ^ message[82] ^ message[83] ^ message[112] ^ message[113] ^ message[114] ^ message[115] ^ message[116] ^ message[117] ^ message[118] ^ message[119] ^ message[176] ^ message[177] ^ message[178] ^ message[179] ^ message[180] ^ message[181] ^ message[182] ^ message[183] ^ message[184] ^ message[185] ^ message[186] ^ message[187] ^ message[188] ^ message[189] ^ message[190] ^ message[191] ^ message[192] ^ message[193] ^ message[194] ^ message[195] ^ message[196] ^ message[197] ^ message[198] ^ message[199] ^ message[200] ^ message[201] ^ message[202] ^ message[203] ^ message[204] ^ message[205] ^ message[206] ^ message[207] ^ message[208] ^ message[209] ^ message[210] ^ message[211] ^ message[212] ^ message[213] ^ message[214] ^ message[215] ^ message[216] ^ message[217] ^ message[218] ^ message[219] ^ message[220] ^ message[221] ^ message[222] ^ message[223] ^ message[224] ^ message[225] ^ message[226] ^ message[227] ^ message[228] ^ message[229] ^ message[230] ^ message[231] ^ message[232] ^ message[233] ^ message[234] ^ message[235] ^ message[236] ^ message[237] ^ message[238] ^ message[239] ^ message[240] ^ message[241] ^ message[242] ^ message[243] ^ message[244] ^ message[245];
    assign parity[2] = message[35] ^ message[36] ^ message[37] ^ message[38] ^ message[39] ^ message[40] ^ message[41] ^ message[42] ^ message[43] ^ message[44] ^ message[45] ^ message[46] ^ message[47] ^ message[48] ^ message[49] ^ message[50] ^ message[51] ^ message[52] ^ message[53] ^ message[54] ^ message[55] ^ message[77] ^ message[78] ^ message[79] ^ message[80] ^ message[81] ^ message[82] ^ message[83] ^ message[105] ^ message[106] ^ message[107] ^ message[108] ^ message[109] ^ message[110] ^ message[111] ^ message[119] ^ message[141] ^ message[142] ^ message[143] ^ message[144] ^ message[145] ^ message[146] ^ message[147] ^ message[148] ^ message[149] ^ message[150] ^ message[151] ^ message[152] ^ message[153] ^ message[154] ^ message[155] ^ message[156] ^ message[157] ^ message[158] ^ message[159] ^ message[160] ^ message[161] ^ message[162] ^ message[163] ^ message[164] ^ message[165] ^ message[166] ^ message[167] ^ message[168] ^ message[169] ^ message[170] ^ message[171] ^ message[172] ^ message[173] ^ message[174] ^ message[175] ^ message[211] ^ message[212] ^ message[213] ^ message[214] ^ message[215] ^ message[216] ^ message[217] ^ message[218] ^ message[219] ^ message[220] ^ message[221] ^ message[222] ^ message[223] ^ message[224] ^ message[225] ^ message[226] ^ message[227] ^ message[228] ^ message[229] ^ message[230] ^ message[231] ^ message[232] ^ message[233] ^ message[234] ^ message[235] ^ message[236] ^ message[237] ^ message[238] ^ message[239] ^ message[240] ^ message[241] ^ message[242] ^ message[243] ^ message[244] ^ message[245];
    assign parity[3] = message[20] ^ message[21] ^ message[22] ^ message[23] ^ message[24] ^ message[25] ^ message[26] ^ message[27] ^ message[28] ^ message[29] ^ message[30] ^ message[31] ^ message[32] ^ message[33] ^ message[34] ^ message[50] ^ message[51] ^ message[52] ^ message[53] ^ message[54] ^ message[55] ^ message[71] ^ message[72] ^ message[73] ^ message[74] ^ message[75] ^ message[76] ^ message[83] ^ message[99] ^ message[100] ^ message[101] ^ message[102] ^ message[103] ^ message[104] ^ message[111] ^ message[118] ^ message[126] ^ message[127] ^ message[128] ^ message[129] ^ message[130] ^ message[131] ^ message[132] ^ message[133] ^ message[134] ^ message[135] ^ message[136] ^ message[137] ^ message[138] ^ message[139] ^ message[140] ^ message[156] ^ message[157] ^ message[158] ^ message[159] ^ message[160] ^ message[161] ^ message[162] ^ message[163] ^ message[164] ^ message[165] ^ message[166] ^ message[167] ^ message[168] ^ message[169] ^ message[170] ^ message[171] ^ message[172] ^ message[173] ^ message[174] ^ message[175] ^ message[191] ^ message[192] ^ message[193] ^ message[194] ^ message[195] ^ message[196] ^ message[197] ^ message[198] ^ message[199] ^ message[200] ^ message[201] ^ message[202] ^ message[203] ^ message[204] ^ message[205] ^ message[206] ^ message[207] ^ message[208] ^ message[209] ^ message[210] ^ message[231] ^ message[232] ^ message[233] ^ message[234] ^ message[235] ^ message[236] ^ message[237] ^ message[238] ^ message[239] ^ message[240] ^ message[241] ^ message[242] ^ message[243] ^ message[244] ^ message[245];
    assign parity[4] = message[10] ^ message[11] ^ message[12] ^ message[13] ^ message[14] ^ message[15] ^ message[16] ^ message[17] ^ message[18] ^ message[19] ^ message[30] ^ message[31] ^ message[32] ^ message[33] ^ message[34] ^ message[45] ^ message[46] ^ message[47] ^ message[48] ^ message[49] ^ message[55] ^ message[66] ^ message[67] ^ message[68] ^ message[69] ^ message[70] ^ message[76] ^ message[82] ^ message[94] ^ message[95] ^ message[96] ^ message[97] ^ message[98] ^ message[104] ^ message[110] ^ message[117] ^ message[121] ^ message[122] ^ message[123] ^ message[124] ^ message[125] ^ message[131] ^ message[132] ^ message[133] ^ message[134] ^ message[135] ^ message[136] ^ message[137] ^ message[138] ^ message[139] ^ message[140] ^ message[146] ^ message[147] ^ message[148] ^ message[149] ^ message[150] ^ message[151] ^ message[152] ^ message[153] ^ message[154] ^ message[155] ^ message[166] ^ message[167] ^ message[168] ^ message[169] ^ message[170] ^ message[171] ^ message[172] ^ message[173] ^ message[174] ^ message[175] ^ message[181] ^ message[182] ^ message[183] ^ message[184] ^ message[185] ^ message[186] ^ message[187] ^ message[188] ^ message[189] ^ message[190] ^ message[201] ^ message[202] ^ message[203] ^ message[204] ^ message[205] ^ message[206] ^ message[207] ^ message[208] ^ message[209] ^ message[210] ^ message[221] ^ message[222] ^ message[223] ^ message[224] ^ message[225] ^ message[226] ^ message[227] ^ message[228] ^ message[229] ^ message[230] ^ message[241] ^ message[242] ^ message[243] ^ message[244] ^ message[245] ^ message[251] ^ message[252] ^ message[253] ^ message[254] ^ message[255];
    assign parity[5] = message[4] ^ message[5] ^ message[6] ^ message[7] ^ message[8] ^ message[9] ^ message[16] ^ message[17] ^ message[18] ^ message[19] ^ message[26] ^ message[27] ^ message[28] ^ message[29] ^ message[34] ^ message[41] ^ message[42] ^ message[43] ^ message[44] ^ message[49] ^ message[54] ^ message[62] ^ message[63] ^ message[64] ^ message[65] ^ message[70] ^ message[75] ^ message[81] ^ message[90] ^ message[91] ^ message[92] ^ message[93] ^ message[98] ^ message[103] ^ message[109] ^ message[116] ^ message[120] ^ message[122] ^ message[123] ^ message[124] ^ message[125] ^ message[127] ^ message[128] ^ message[129] ^ message[130] ^ message[135] ^ message[136] ^ message[137] ^ message[138] ^ message[139] ^ message[140] ^ message[142] ^ message[143] ^ message[144] ^ message[145] ^ message[150] ^ message[151] ^ message[152] ^ message[153] ^ message[154] ^ message[155] ^ message[160] ^ message[161] ^ message[162] ^ message[163] ^ message[164] ^ message[165] ^ message[172] ^ message[173] ^ message[174] ^ message[175] ^ message[177] ^ message[178] ^ message[179] ^ message[180] ^ message[185] ^ message[186] ^ message[187] ^ message[188] ^ message[189] ^ message[190] ^ message[195] ^ message[196] ^ message[197] ^ message[198] ^ message[199] ^ message[200] ^ message[207] ^ message[208] ^ message[209] ^ message[210] ^ message[215] ^ message[216] ^ message[217] ^ message[218] ^ message[219] ^ message[220] ^ message[227] ^ message[228] ^ message[229] ^ message[230] ^ message[237] ^ message[238] ^ message[239] ^ message[240] ^ message[245] ^ message[247] ^ message[248] ^ message[249] ^ message[250] ^ message[255];
    assign parity[6] = message[1] ^ message[2] ^ message[3] ^ message[7] ^ message[8] ^ message[9] ^ message[13] ^ message[14] ^ message[15] ^ message[19] ^ message[23] ^ message[24] ^ message[25] ^ message[29] ^ message[33] ^ message[38] ^ message[39] ^ message[40] ^ message[44] ^ message[48] ^ message[53] ^ message[59] ^ message[60] ^ message[61] ^ message[65] ^ message[69] ^ message[74] ^ message[80] ^ message[87] ^ message[88] ^ message[89] ^ message[93] ^ message[97] ^ message[102] ^ message[108] ^ message[115] ^ message[120] ^ message[121] ^ message[123] ^ message[124] ^ message[125] ^ message[126] ^ message[128] ^ message[129] ^ message[130] ^ message[132] ^ message[133] ^ message[134] ^ message[138] ^ message[139] ^ message[140] ^ message[141] ^ message[143] ^ message[144] ^ message[145] ^ message[147] ^ message[148] ^ message[149] ^ message[153] ^ message[154] ^ message[155] ^ message[157] ^ message[158] ^ message[159] ^ message[163] ^ message[164] ^ message[165] ^ message[169] ^ message[170] ^ message[171] ^ message[175] ^ message[176] ^ message[178] ^ message[179] ^ message[180] ^ message[182] ^ message[183] ^ message[184] ^ message[188] ^ message[189] ^ message[190] ^ message[192] ^ message[193] ^ message[194] ^ message[198] ^ message[199] ^ message[200] ^ message[204] ^ message[205] ^ message[206] ^ message[210] ^ message[212] ^ message[213] ^ message[214] ^ message[218] ^ message[219] ^ message[220] ^ message[224] ^ message[225] ^ message[226] ^ message[230] ^ message[234] ^ message[235] ^ message[236] ^ message[240] ^ message[244] ^ message[246] ^ message[248] ^ message[249] ^ message[250] ^ message[252] ^ message[253] ^ message[254];
    assign parity[7] = message[0] ^ message[2] ^ message[3] ^ message[5] ^ message[6] ^ message[9] ^ message[11] ^ message[12] ^ message[15] ^ message[18] ^ message[21] ^ message[22] ^ message[25] ^ message[28] ^ message[32] ^ message[36] ^ message[37] ^ message[40] ^ message[43] ^ message[47] ^ message[52] ^ message[57] ^ message[58] ^ message[61] ^ message[64] ^ message[68] ^ message[73] ^ message[79] ^ message[85] ^ message[86] ^ message[89] ^ message[92] ^ message[96] ^ message[101] ^ message[107] ^ message[114] ^ message[120] ^ message[121] ^ message[122] ^ message[124] ^ message[125] ^ message[126] ^ message[127] ^ message[129] ^ message[130] ^ message[131] ^ message[133] ^ message[134] ^ message[136] ^ message[137] ^ message[140] ^ message[141] ^ message[142] ^ message[144] ^ message[145] ^ message[146] ^ message[148] ^ message[149] ^ message[151] ^ message[152] ^ message[155] ^ message[156] ^ message[158] ^ message[159] ^ message[161] ^ message[162] ^ message[165] ^ message[167] ^ message[168] ^ message[171] ^ message[174] ^ message[176] ^ message[177] ^ message[179] ^ message[180] ^ message[181] ^ message[183] ^ message[184] ^ message[186] ^ message[187] ^ message[190] ^ message[191] ^ message[193] ^ message[194] ^ message[196] ^ message[197] ^ message[200] ^ message[202] ^ message[203] ^ message[206] ^ message[209] ^ message[211] ^ message[213] ^ message[214] ^ message[216] ^ message[217] ^ message[220] ^ message[222] ^ message[223] ^ message[226] ^ message[229] ^ message[232] ^ message[233] ^ message[236] ^ message[239] ^ message[243] ^ message[246] ^ message[247] ^ message[249] ^ message[250] ^ message[251] ^ message[253] ^ message[254];
    assign parity[8] = message[0] ^ message[1] ^ message[3] ^ message[4] ^ message[6] ^ message[8] ^ message[10] ^ message[12] ^ message[14] ^ message[17] ^ message[20] ^ message[22] ^ message[24] ^ message[27] ^ message[31] ^ message[35] ^ message[37] ^ message[39] ^ message[42] ^ message[46] ^ message[51] ^ message[56] ^ message[58] ^ message[60] ^ message[63] ^ message[67] ^ message[72] ^ message[78] ^ message[84] ^ message[86] ^ message[88] ^ message[91] ^ message[95] ^ message[100] ^ message[106] ^ message[113] ^ message[120] ^ message[121] ^ message[122] ^ message[123] ^ message[125] ^ message[126] ^ message[127] ^ message[128] ^ message[130] ^ message[131] ^ message[132] ^ message[134] ^ message[135] ^ message[137] ^ message[139] ^ message[141] ^ message[142] ^ message[143] ^ message[145] ^ message[146] ^ message[147] ^ message[149] ^ message[150] ^ message[152] ^ message[154] ^ message[156] ^ message[157] ^ message[159] ^ message[160] ^ message[162] ^ message[164] ^ message[166] ^ message[168] ^ message[170] ^ message[173] ^ message[176] ^ message[177] ^ message[178] ^ message[180] ^ message[181] ^ message[182] ^ message[184] ^ message[185] ^ message[187] ^ message[189] ^ message[191] ^ message[192] ^ message[194] ^ message[195] ^ message[197] ^ message[199] ^ message[201] ^ message[203] ^ message[205] ^ message[208] ^ message[211] ^ message[212] ^ message[214] ^ message[215] ^ message[217] ^ message[219] ^ message[221] ^ message[223] ^ message[225] ^ message[228] ^ message[231] ^ message[233] ^ message[235] ^ message[238] ^ message[242] ^ message[246] ^ message[247] ^ message[248] ^ message[250] ^ message[251] ^ message[252] ^ message[254] ^ message[255];
    assign parity[9] = message[0] ^ message[1] ^ message[2] ^ message[4] ^ message[5] ^ message[7] ^ message[10] ^ message[11] ^ message[13] ^ message[16] ^ message[20] ^ message[21] ^ message[23] ^ message[26] ^ message[30] ^ message[35] ^ message[36] ^ message[38] ^ message[41] ^ message[45] ^ message[50] ^ message[56] ^ message[57] ^ message[59] ^ message[62] ^ message[66] ^ message[71] ^ message[77] ^ message[84] ^ message[85] ^ message[87] ^ message[90] ^ message[94] ^ message[99] ^ message[105] ^ message[112] ^ message[120] ^ message[121] ^ message[122] ^ message[123] ^ message[124] ^ message[126] ^ message[127] ^ message[128] ^ message[129] ^ message[131] ^ message[132] ^ message[133] ^ message[135] ^ message[136] ^ message[138] ^ message[141] ^ message[142] ^ message[143] ^ message[144] ^ message[146] ^ message[147] ^ message[148] ^ message[150] ^ message[151] ^ message[153] ^ message[156] ^ message[157] ^ message[158] ^ message[160] ^ message[161] ^ message[163] ^ message[166] ^ message[167] ^ message[169] ^ message[172] ^ message[176] ^ message[177] ^ message[178] ^ message[179] ^ message[181] ^ message[182] ^ message[183] ^ message[185] ^ message[186] ^ message[188] ^ message[191] ^ message[192] ^ message[193] ^ message[195] ^ message[196] ^ message[198] ^ message[201] ^ message[202] ^ message[204] ^ message[207] ^ message[211] ^ message[212] ^ message[213] ^ message[215] ^ message[216] ^ message[218] ^ message[221] ^ message[222] ^ message[224] ^ message[227] ^ message[231] ^ message[232] ^ message[234] ^ message[237] ^ message[241] ^ message[246] ^ message[247] ^ message[248] ^ message[249] ^ message[251] ^ message[252] ^ message[253] ^ message[255];
  end else if ((CodewordWidth == 523) && (MessageWidth == 512)) begin : gen_523_512
    `BR_ASSERT_STATIC(parity_width_matches_a, ParityWidth == 11)
    assign parity[0] = message[120] ^ message[121] ^ message[122] ^ message[123] ^ message[124] ^ message[125] ^ message[126] ^ message[127] ^ message[128] ^ message[129] ^ message[130] ^ message[131] ^ message[132] ^ message[133] ^ message[134] ^ message[135] ^ message[136] ^ message[137] ^ message[138] ^ message[139] ^ message[140] ^ message[141] ^ message[142] ^ message[143] ^ message[144] ^ message[145] ^ message[146] ^ message[147] ^ message[148] ^ message[149] ^ message[150] ^ message[151] ^ message[152] ^ message[153] ^ message[154] ^ message[155] ^ message[156] ^ message[157] ^ message[158] ^ message[159] ^ message[160] ^ message[161] ^ message[162] ^ message[163] ^ message[164] ^ message[417] ^ message[418] ^ message[419] ^ message[420] ^ message[421] ^ message[422] ^ message[423] ^ message[424] ^ message[425] ^ message[426] ^ message[427] ^ message[428] ^ message[429] ^ message[430] ^ message[431] ^ message[432] ^ message[433] ^ message[434] ^ message[435] ^ message[436] ^ message[437] ^ message[438] ^ message[439] ^ message[440] ^ message[441] ^ message[442] ^ message[443] ^ message[444] ^ message[445] ^ message[446] ^ message[447] ^ message[448] ^ message[449] ^ message[450] ^ message[451] ^ message[452] ^ message[453] ^ message[454] ^ message[455] ^ message[456] ^ message[457] ^ message[458] ^ message[459] ^ message[460] ^ message[461] ^ message[462] ^ message[463] ^ message[464] ^ message[465] ^ message[466] ^ message[467] ^ message[468] ^ message[469] ^ message[470] ^ message[471] ^ message[472] ^ message[473] ^ message[474] ^ message[475] ^ message[476] ^ message[477] ^ message[478] ^ message[479] ^ message[480] ^ message[481] ^ message[482] ^ message[483] ^ message[484] ^ message[485] ^ message[486] ^ message[487] ^ message[488] ^ message[489] ^ message[490] ^ message[491] ^ message[492] ^ message[493] ^ message[494] ^ message[495] ^ message[496] ^ message[497] ^ message[498] ^ message[499] ^ message[500] ^ message[501] ^ message[502] ^ message[503] ^ message[504] ^ message[505] ^ message[506] ^ message[507] ^ message[508] ^ message[509] ^ message[510] ^ message[511];
    assign parity[1] = message[84] ^ message[85] ^ message[86] ^ message[87] ^ message[88] ^ message[89] ^ message[90] ^ message[91] ^ message[92] ^ message[93] ^ message[94] ^ message[95] ^ message[96] ^ message[97] ^ message[98] ^ message[99] ^ message[100] ^ message[101] ^ message[102] ^ message[103] ^ message[104] ^ message[105] ^ message[106] ^ message[107] ^ message[108] ^ message[109] ^ message[110] ^ message[111] ^ message[112] ^ message[113] ^ message[114] ^ message[115] ^ message[116] ^ message[117] ^ message[118] ^ message[119] ^ message[156] ^ message[157] ^ message[158] ^ message[159] ^ message[160] ^ message[161] ^ message[162] ^ message[163] ^ message[164] ^ message[291] ^ message[292] ^ message[293] ^ message[294] ^ message[295] ^ message[296] ^ message[297] ^ message[298] ^ message[299] ^ message[300] ^ message[301] ^ message[302] ^ message[303] ^ message[304] ^ message[305] ^ message[306] ^ message[307] ^ message[308] ^ message[309] ^ message[310] ^ message[311] ^ message[312] ^ message[313] ^ message[314] ^ message[315] ^ message[316] ^ message[317] ^ message[318] ^ message[319] ^ message[320] ^ message[321] ^ message[322] ^ message[323] ^ message[324] ^ message[325] ^ message[326] ^ message[327] ^ message[328] ^ message[329] ^ message[330] ^ message[331] ^ message[332] ^ message[333] ^ message[334] ^ message[335] ^ message[336] ^ message[337] ^ message[338] ^ message[339] ^ message[340] ^ message[341] ^ message[342] ^ message[343] ^ message[344] ^ message[345] ^ message[346] ^ message[347] ^ message[348] ^ message[349] ^ message[350] ^ message[351] ^ message[352] ^ message[353] ^ message[354] ^ message[355] ^ message[356] ^ message[357] ^ message[358] ^ message[359] ^ message[360] ^ message[361] ^ message[362] ^ message[363] ^ message[364] ^ message[365] ^ message[366] ^ message[367] ^ message[368] ^ message[369] ^ message[370] ^ message[371] ^ message[372] ^ message[373] ^ message[374] ^ message[375] ^ message[376] ^ message[377] ^ message[378] ^ message[379] ^ message[380] ^ message[381] ^ message[382] ^ message[383] ^ message[384] ^ message[385] ^ message[386] ^ message[387] ^ message[388] ^ message[389] ^ message[390] ^ message[391] ^ message[392] ^ message[393] ^ message[394] ^ message[395] ^ message[396] ^ message[397] ^ message[398] ^ message[399] ^ message[400] ^ message[401] ^ message[402] ^ message[403] ^ message[404] ^ message[405] ^ message[406] ^ message[407] ^ message[408] ^ message[409] ^ message[410] ^ message[411] ^ message[412] ^ message[413] ^ message[414] ^ message[415] ^ message[416];
    assign parity[2] = message[56] ^ message[57] ^ message[58] ^ message[59] ^ message[60] ^ message[61] ^ message[62] ^ message[63] ^ message[64] ^ message[65] ^ message[66] ^ message[67] ^ message[68] ^ message[69] ^ message[70] ^ message[71] ^ message[72] ^ message[73] ^ message[74] ^ message[75] ^ message[76] ^ message[77] ^ message[78] ^ message[79] ^ message[80] ^ message[81] ^ message[82] ^ message[83] ^ message[112] ^ message[113] ^ message[114] ^ message[115] ^ message[116] ^ message[117] ^ message[118] ^ message[119] ^ message[148] ^ message[149] ^ message[150] ^ message[151] ^ message[152] ^ message[153] ^ message[154] ^ message[155] ^ message[164] ^ message[221] ^ message[222] ^ message[223] ^ message[224] ^ message[225] ^ message[226] ^ message[227] ^ message[228] ^ message[229] ^ message[230] ^ message[231] ^ message[232] ^ message[233] ^ message[234] ^ message[235] ^ message[236] ^ message[237] ^ message[238] ^ message[239] ^ message[240] ^ message[241] ^ message[242] ^ message[243] ^ message[244] ^ message[245] ^ message[246] ^ message[247] ^ message[248] ^ message[249] ^ message[250] ^ message[251] ^ message[252] ^ message[253] ^ message[254] ^ message[255] ^ message[256] ^ message[257] ^ message[258] ^ message[259] ^ message[260] ^ message[261] ^ message[262] ^ message[263] ^ message[264] ^ message[265] ^ message[266] ^ message[267] ^ message[268] ^ message[269] ^ message[270] ^ message[271] ^ message[272] ^ message[273] ^ message[274] ^ message[275] ^ message[276] ^ message[277] ^ message[278] ^ message[279] ^ message[280] ^ message[281] ^ message[282] ^ message[283] ^ message[284] ^ message[285] ^ message[286] ^ message[287] ^ message[288] ^ message[289] ^ message[290] ^ message[361] ^ message[362] ^ message[363] ^ message[364] ^ message[365] ^ message[366] ^ message[367] ^ message[368] ^ message[369] ^ message[370] ^ message[371] ^ message[372] ^ message[373] ^ message[374] ^ message[375] ^ message[376] ^ message[377] ^ message[378] ^ message[379] ^ message[380] ^ message[381] ^ message[382] ^ message[383] ^ message[384] ^ message[385] ^ message[386] ^ message[387] ^ message[388] ^ message[389] ^ message[390] ^ message[391] ^ message[392] ^ message[393] ^ message[394] ^ message[395] ^ message[396] ^ message[397] ^ message[398] ^ message[399] ^ message[400] ^ message[401] ^ message[402] ^ message[403] ^ message[404] ^ message[405] ^ message[406] ^ message[407] ^ message[408] ^ message[409] ^ message[410] ^ message[411] ^ message[412] ^ message[413] ^ message[414] ^ message[415] ^ message[416] ^ message[487] ^ message[488] ^ message[489] ^ message[490] ^ message[491] ^ message[492] ^ message[493] ^ message[494] ^ message[495] ^ message[496] ^ message[497] ^ message[498] ^ message[499] ^ message[500] ^ message[501] ^ message[502] ^ message[503] ^ message[504] ^ message[505] ^ message[506] ^ message[507] ^ message[508] ^ message[509] ^ message[510] ^ message[511];
    assign parity[3] = message[35] ^ message[36] ^ message[37] ^ message[38] ^ message[39] ^ message[40] ^ message[41] ^ message[42] ^ message[43] ^ message[44] ^ message[45] ^ message[46] ^ message[47] ^ message[48] ^ message[49] ^ message[50] ^ message[51] ^ message[52] ^ message[53] ^ message[54] ^ message[55] ^ message[77] ^ message[78] ^ message[79] ^ message[80] ^ message[81] ^ message[82] ^ message[83] ^ message[105] ^ message[106] ^ message[107] ^ message[108] ^ message[109] ^ message[110] ^ message[111] ^ message[119] ^ message[141] ^ message[142] ^ message[143] ^ message[144] ^ message[145] ^ message[146] ^ message[147] ^ message[155] ^ message[163] ^ message[186] ^ message[187] ^ message[188] ^ message[189] ^ message[190] ^ message[191] ^ message[192] ^ message[193] ^ message[194] ^ message[195] ^ message[196] ^ message[197] ^ message[198] ^ message[199] ^ message[200] ^ message[201] ^ message[202] ^ message[203] ^ message[204] ^ message[205] ^ message[206] ^ message[207] ^ message[208] ^ message[209] ^ message[210] ^ message[211] ^ message[212] ^ message[213] ^ message[214] ^ message[215] ^ message[216] ^ message[217] ^ message[218] ^ message[219] ^ message[220] ^ message[256] ^ message[257] ^ message[258] ^ message[259] ^ message[260] ^ message[261] ^ message[262] ^ message[263] ^ message[264] ^ message[265] ^ message[266] ^ message[267] ^ message[268] ^ message[269] ^ message[270] ^ message[271] ^ message[272] ^ message[273] ^ message[274] ^ message[275] ^ message[276] ^ message[277] ^ message[278] ^ message[279] ^ message[280] ^ message[281] ^ message[282] ^ message[283] ^ message[284] ^ message[285] ^ message[286] ^ message[287] ^ message[288] ^ message[289] ^ message[290] ^ message[326] ^ message[327] ^ message[328] ^ message[329] ^ message[330] ^ message[331] ^ message[332] ^ message[333] ^ message[334] ^ message[335] ^ message[336] ^ message[337] ^ message[338] ^ message[339] ^ message[340] ^ message[341] ^ message[342] ^ message[343] ^ message[344] ^ message[345] ^ message[346] ^ message[347] ^ message[348] ^ message[349] ^ message[350] ^ message[351] ^ message[352] ^ message[353] ^ message[354] ^ message[355] ^ message[356] ^ message[357] ^ message[358] ^ message[359] ^ message[360] ^ message[396] ^ message[397] ^ message[398] ^ message[399] ^ message[400] ^ message[401] ^ message[402] ^ message[403] ^ message[404] ^ message[405] ^ message[406] ^ message[407] ^ message[408] ^ message[409] ^ message[410] ^ message[411] ^ message[412] ^ message[413] ^ message[414] ^ message[415] ^ message[416] ^ message[452] ^ message[453] ^ message[454] ^ message[455] ^ message[456] ^ message[457] ^ message[458] ^ message[459] ^ message[460] ^ message[461] ^ message[462] ^ message[463] ^ message[464] ^ message[465] ^ message[466] ^ message[467] ^ message[468] ^ message[469] ^ message[470] ^ message[471] ^ message[472] ^ message[473] ^ message[474] ^ message[475] ^ message[476] ^ message[477] ^ message[478] ^ message[479] ^ message[480] ^ message[481] ^ message[482] ^ message[483] ^ message[484] ^ message[485] ^ message[486];
    assign parity[4] = message[20] ^ message[21] ^ message[22] ^ message[23] ^ message[24] ^ message[25] ^ message[26] ^ message[27] ^ message[28] ^ message[29] ^ message[30] ^ message[31] ^ message[32] ^ message[33] ^ message[34] ^ message[50] ^ message[51] ^ message[52] ^ message[53] ^ message[54] ^ message[55] ^ message[71] ^ message[72] ^ message[73] ^ message[74] ^ message[75] ^ message[76] ^ message[83] ^ message[99] ^ message[100] ^ message[101] ^ message[102] ^ message[103] ^ message[104] ^ message[111] ^ message[118] ^ message[135] ^ message[136] ^ message[137] ^ message[138] ^ message[139] ^ message[140] ^ message[147] ^ message[154] ^ message[162] ^ message[171] ^ message[172] ^ message[173] ^ message[174] ^ message[175] ^ message[176] ^ message[177] ^ message[178] ^ message[179] ^ message[180] ^ message[181] ^ message[182] ^ message[183] ^ message[184] ^ message[185] ^ message[201] ^ message[202] ^ message[203] ^ message[204] ^ message[205] ^ message[206] ^ message[207] ^ message[208] ^ message[209] ^ message[210] ^ message[211] ^ message[212] ^ message[213] ^ message[214] ^ message[215] ^ message[216] ^ message[217] ^ message[218] ^ message[219] ^ message[220] ^ message[236] ^ message[237] ^ message[238] ^ message[239] ^ message[240] ^ message[241] ^ message[242] ^ message[243] ^ message[244] ^ message[245] ^ message[246] ^ message[247] ^ message[248] ^ message[249] ^ message[250] ^ message[251] ^ message[252] ^ message[253] ^ message[254] ^ message[255] ^ message[276] ^ message[277] ^ message[278] ^ message[279] ^ message[280] ^ message[281] ^ message[282] ^ message[283] ^ message[284] ^ message[285] ^ message[286] ^ message[287] ^ message[288] ^ message[289] ^ message[290] ^ message[306] ^ message[307] ^ message[308] ^ message[309] ^ message[310] ^ message[311] ^ message[312] ^ message[313] ^ message[314] ^ message[315] ^ message[316] ^ message[317] ^ message[318] ^ message[319] ^ message[320] ^ message[321] ^ message[322] ^ message[323] ^ message[324] ^ message[325] ^ message[346] ^ message[347] ^ message[348] ^ message[349] ^ message[350] ^ message[351] ^ message[352] ^ message[353] ^ message[354] ^ message[355] ^ message[356] ^ message[357] ^ message[358] ^ message[359] ^ message[360] ^ message[381] ^ message[382] ^ message[383] ^ message[384] ^ message[385] ^ message[386] ^ message[387] ^ message[388] ^ message[389] ^ message[390] ^ message[391] ^ message[392] ^ message[393] ^ message[394] ^ message[395] ^ message[411] ^ message[412] ^ message[413] ^ message[414] ^ message[415] ^ message[416] ^ message[432] ^ message[433] ^ message[434] ^ message[435] ^ message[436] ^ message[437] ^ message[438] ^ message[439] ^ message[440] ^ message[441] ^ message[442] ^ message[443] ^ message[444] ^ message[445] ^ message[446] ^ message[447] ^ message[448] ^ message[449] ^ message[450] ^ message[451] ^ message[472] ^ message[473] ^ message[474] ^ message[475] ^ message[476] ^ message[477] ^ message[478] ^ message[479] ^ message[480] ^ message[481] ^ message[482] ^ message[483] ^ message[484] ^ message[485] ^ message[486] ^ message[507] ^ message[508] ^ message[509] ^ message[510] ^ message[511];
    assign parity[5] = message[10] ^ message[11] ^ message[12] ^ message[13] ^ message[14] ^ message[15] ^ message[16] ^ message[17] ^ message[18] ^ message[19] ^ message[30] ^ message[31] ^ message[32] ^ message[33] ^ message[34] ^ message[45] ^ message[46] ^ message[47] ^ message[48] ^ message[49] ^ message[55] ^ message[66] ^ message[67] ^ message[68] ^ message[69] ^ message[70] ^ message[76] ^ message[82] ^ message[94] ^ message[95] ^ message[96] ^ message[97] ^ message[98] ^ message[104] ^ message[110] ^ message[117] ^ message[130] ^ message[131] ^ message[132] ^ message[133] ^ message[134] ^ message[140] ^ message[146] ^ message[153] ^ message[161] ^ message[166] ^ message[167] ^ message[168] ^ message[169] ^ message[170] ^ message[176] ^ message[177] ^ message[178] ^ message[179] ^ message[180] ^ message[181] ^ message[182] ^ message[183] ^ message[184] ^ message[185] ^ message[191] ^ message[192] ^ message[193] ^ message[194] ^ message[195] ^ message[196] ^ message[197] ^ message[198] ^ message[199] ^ message[200] ^ message[211] ^ message[212] ^ message[213] ^ message[214] ^ message[215] ^ message[216] ^ message[217] ^ message[218] ^ message[219] ^ message[220] ^ message[226] ^ message[227] ^ message[228] ^ message[229] ^ message[230] ^ message[231] ^ message[232] ^ message[233] ^ message[234] ^ message[235] ^ message[246] ^ message[247] ^ message[248] ^ message[249] ^ message[250] ^ message[251] ^ message[252] ^ message[253] ^ message[254] ^ message[255] ^ message[266] ^ message[267] ^ message[268] ^ message[269] ^ message[270] ^ message[271] ^ message[272] ^ message[273] ^ message[274] ^ message[275] ^ message[286] ^ message[287] ^ message[288] ^ message[289] ^ message[290] ^ message[296] ^ message[297] ^ message[298] ^ message[299] ^ message[300] ^ message[301] ^ message[302] ^ message[303] ^ message[304] ^ message[305] ^ message[316] ^ message[317] ^ message[318] ^ message[319] ^ message[320] ^ message[321] ^ message[322] ^ message[323] ^ message[324] ^ message[325] ^ message[336] ^ message[337] ^ message[338] ^ message[339] ^ message[340] ^ message[341] ^ message[342] ^ message[343] ^ message[344] ^ message[345] ^ message[356] ^ message[357] ^ message[358] ^ message[359] ^ message[360] ^ message[371] ^ message[372] ^ message[373] ^ message[374] ^ message[375] ^ message[376] ^ message[377] ^ message[378] ^ message[379] ^ message[380] ^ message[391] ^ message[392] ^ message[393] ^ message[394] ^ message[395] ^ message[406] ^ message[407] ^ message[408] ^ message[409] ^ message[410] ^ message[416] ^ message[422] ^ message[423] ^ message[424] ^ message[425] ^ message[426] ^ message[427] ^ message[428] ^ message[429] ^ message[430] ^ message[431] ^ message[442] ^ message[443] ^ message[444] ^ message[445] ^ message[446] ^ message[447] ^ message[448] ^ message[449] ^ message[450] ^ message[451] ^ message[462] ^ message[463] ^ message[464] ^ message[465] ^ message[466] ^ message[467] ^ message[468] ^ message[469] ^ message[470] ^ message[471] ^ message[482] ^ message[483] ^ message[484] ^ message[485] ^ message[486] ^ message[497] ^ message[498] ^ message[499] ^ message[500] ^ message[501] ^ message[502] ^ message[503] ^ message[504] ^ message[505] ^ message[506];
    assign parity[6] = message[4] ^ message[5] ^ message[6] ^ message[7] ^ message[8] ^ message[9] ^ message[16] ^ message[17] ^ message[18] ^ message[19] ^ message[26] ^ message[27] ^ message[28] ^ message[29] ^ message[34] ^ message[41] ^ message[42] ^ message[43] ^ message[44] ^ message[49] ^ message[54] ^ message[62] ^ message[63] ^ message[64] ^ message[65] ^ message[70] ^ message[75] ^ message[81] ^ message[90] ^ message[91] ^ message[92] ^ message[93] ^ message[98] ^ message[103] ^ message[109] ^ message[116] ^ message[126] ^ message[127] ^ message[128] ^ message[129] ^ message[134] ^ message[139] ^ message[145] ^ message[152] ^ message[160] ^ message[165] ^ message[167] ^ message[168] ^ message[169] ^ message[170] ^ message[172] ^ message[173] ^ message[174] ^ message[175] ^ message[180] ^ message[181] ^ message[182] ^ message[183] ^ message[184] ^ message[185] ^ message[187] ^ message[188] ^ message[189] ^ message[190] ^ message[195] ^ message[196] ^ message[197] ^ message[198] ^ message[199] ^ message[200] ^ message[205] ^ message[206] ^ message[207] ^ message[208] ^ message[209] ^ message[210] ^ message[217] ^ message[218] ^ message[219] ^ message[220] ^ message[222] ^ message[223] ^ message[224] ^ message[225] ^ message[230] ^ message[231] ^ message[232] ^ message[233] ^ message[234] ^ message[235] ^ message[240] ^ message[241] ^ message[242] ^ message[243] ^ message[244] ^ message[245] ^ message[252] ^ message[253] ^ message[254] ^ message[255] ^ message[260] ^ message[261] ^ message[262] ^ message[263] ^ message[264] ^ message[265] ^ message[272] ^ message[273] ^ message[274] ^ message[275] ^ message[282] ^ message[283] ^ message[284] ^ message[285] ^ message[290] ^ message[292] ^ message[293] ^ message[294] ^ message[295] ^ message[300] ^ message[301] ^ message[302] ^ message[303] ^ message[304] ^ message[305] ^ message[310] ^ message[311] ^ message[312] ^ message[313] ^ message[314] ^ message[315] ^ message[322] ^ message[323] ^ message[324] ^ message[325] ^ message[330] ^ message[331] ^ message[332] ^ message[333] ^ message[334] ^ message[335] ^ message[342] ^ message[343] ^ message[344] ^ message[345] ^ message[352] ^ message[353] ^ message[354] ^ message[355] ^ message[360] ^ message[365] ^ message[366] ^ message[367] ^ message[368] ^ message[369] ^ message[370] ^ message[377] ^ message[378] ^ message[379] ^ message[380] ^ message[387] ^ message[388] ^ message[389] ^ message[390] ^ message[395] ^ message[402] ^ message[403] ^ message[404] ^ message[405] ^ message[410] ^ message[415] ^ message[418] ^ message[419] ^ message[420] ^ message[421] ^ message[426] ^ message[427] ^ message[428] ^ message[429] ^ message[430] ^ message[431] ^ message[436] ^ message[437] ^ message[438] ^ message[439] ^ message[440] ^ message[441] ^ message[448] ^ message[449] ^ message[450] ^ message[451] ^ message[456] ^ message[457] ^ message[458] ^ message[459] ^ message[460] ^ message[461] ^ message[468] ^ message[469] ^ message[470] ^ message[471] ^ message[478] ^ message[479] ^ message[480] ^ message[481] ^ message[486] ^ message[491] ^ message[492] ^ message[493] ^ message[494] ^ message[495] ^ message[496] ^ message[503] ^ message[504] ^ message[505] ^ message[506];
    assign parity[7] = message[1] ^ message[2] ^ message[3] ^ message[7] ^ message[8] ^ message[9] ^ message[13] ^ message[14] ^ message[15] ^ message[19] ^ message[23] ^ message[24] ^ message[25] ^ message[29] ^ message[33] ^ message[38] ^ message[39] ^ message[40] ^ message[44] ^ message[48] ^ message[53] ^ message[59] ^ message[60] ^ message[61] ^ message[65] ^ message[69] ^ message[74] ^ message[80] ^ message[87] ^ message[88] ^ message[89] ^ message[93] ^ message[97] ^ message[102] ^ message[108] ^ message[115] ^ message[123] ^ message[124] ^ message[125] ^ message[129] ^ message[133] ^ message[138] ^ message[144] ^ message[151] ^ message[159] ^ message[165] ^ message[166] ^ message[168] ^ message[169] ^ message[170] ^ message[171] ^ message[173] ^ message[174] ^ message[175] ^ message[177] ^ message[178] ^ message[179] ^ message[183] ^ message[184] ^ message[185] ^ message[186] ^ message[188] ^ message[189] ^ message[190] ^ message[192] ^ message[193] ^ message[194] ^ message[198] ^ message[199] ^ message[200] ^ message[202] ^ message[203] ^ message[204] ^ message[208] ^ message[209] ^ message[210] ^ message[214] ^ message[215] ^ message[216] ^ message[220] ^ message[221] ^ message[223] ^ message[224] ^ message[225] ^ message[227] ^ message[228] ^ message[229] ^ message[233] ^ message[234] ^ message[235] ^ message[237] ^ message[238] ^ message[239] ^ message[243] ^ message[244] ^ message[245] ^ message[249] ^ message[250] ^ message[251] ^ message[255] ^ message[257] ^ message[258] ^ message[259] ^ message[263] ^ message[264] ^ message[265] ^ message[269] ^ message[270] ^ message[271] ^ message[275] ^ message[279] ^ message[280] ^ message[281] ^ message[285] ^ message[289] ^ message[291] ^ message[293] ^ message[294] ^ message[295] ^ message[297] ^ message[298] ^ message[299] ^ message[303] ^ message[304] ^ message[305] ^ message[307] ^ message[308] ^ message[309] ^ message[313] ^ message[314] ^ message[315] ^ message[319] ^ message[320] ^ message[321] ^ message[325] ^ message[327] ^ message[328] ^ message[329] ^ message[333] ^ message[334] ^ message[335] ^ message[339] ^ message[340] ^ message[341] ^ message[345] ^ message[349] ^ message[350] ^ message[351] ^ message[355] ^ message[359] ^ message[362] ^ message[363] ^ message[364] ^ message[368] ^ message[369] ^ message[370] ^ message[374] ^ message[375] ^ message[376] ^ message[380] ^ message[384] ^ message[385] ^ message[386] ^ message[390] ^ message[394] ^ message[399] ^ message[400] ^ message[401] ^ message[405] ^ message[409] ^ message[414] ^ message[417] ^ message[419] ^ message[420] ^ message[421] ^ message[423] ^ message[424] ^ message[425] ^ message[429] ^ message[430] ^ message[431] ^ message[433] ^ message[434] ^ message[435] ^ message[439] ^ message[440] ^ message[441] ^ message[445] ^ message[446] ^ message[447] ^ message[451] ^ message[453] ^ message[454] ^ message[455] ^ message[459] ^ message[460] ^ message[461] ^ message[465] ^ message[466] ^ message[467] ^ message[471] ^ message[475] ^ message[476] ^ message[477] ^ message[481] ^ message[485] ^ message[488] ^ message[489] ^ message[490] ^ message[494] ^ message[495] ^ message[496] ^ message[500] ^ message[501] ^ message[502] ^ message[506] ^ message[510] ^ message[511];
    assign parity[8] = message[0] ^ message[2] ^ message[3] ^ message[5] ^ message[6] ^ message[9] ^ message[11] ^ message[12] ^ message[15] ^ message[18] ^ message[21] ^ message[22] ^ message[25] ^ message[28] ^ message[32] ^ message[36] ^ message[37] ^ message[40] ^ message[43] ^ message[47] ^ message[52] ^ message[57] ^ message[58] ^ message[61] ^ message[64] ^ message[68] ^ message[73] ^ message[79] ^ message[85] ^ message[86] ^ message[89] ^ message[92] ^ message[96] ^ message[101] ^ message[107] ^ message[114] ^ message[121] ^ message[122] ^ message[125] ^ message[128] ^ message[132] ^ message[137] ^ message[143] ^ message[150] ^ message[158] ^ message[165] ^ message[166] ^ message[167] ^ message[169] ^ message[170] ^ message[171] ^ message[172] ^ message[174] ^ message[175] ^ message[176] ^ message[178] ^ message[179] ^ message[181] ^ message[182] ^ message[185] ^ message[186] ^ message[187] ^ message[189] ^ message[190] ^ message[191] ^ message[193] ^ message[194] ^ message[196] ^ message[197] ^ message[200] ^ message[201] ^ message[203] ^ message[204] ^ message[206] ^ message[207] ^ message[210] ^ message[212] ^ message[213] ^ message[216] ^ message[219] ^ message[221] ^ message[222] ^ message[224] ^ message[225] ^ message[226] ^ message[228] ^ message[229] ^ message[231] ^ message[232] ^ message[235] ^ message[236] ^ message[238] ^ message[239] ^ message[241] ^ message[242] ^ message[245] ^ message[247] ^ message[248] ^ message[251] ^ message[254] ^ message[256] ^ message[258] ^ message[259] ^ message[261] ^ message[262] ^ message[265] ^ message[267] ^ message[268] ^ message[271] ^ message[274] ^ message[277] ^ message[278] ^ message[281] ^ message[284] ^ message[288] ^ message[291] ^ message[292] ^ message[294] ^ message[295] ^ message[296] ^ message[298] ^ message[299] ^ message[301] ^ message[302] ^ message[305] ^ message[306] ^ message[308] ^ message[309] ^ message[311] ^ message[312] ^ message[315] ^ message[317] ^ message[318] ^ message[321] ^ message[324] ^ message[326] ^ message[328] ^ message[329] ^ message[331] ^ message[332] ^ message[335] ^ message[337] ^ message[338] ^ message[341] ^ message[344] ^ message[347] ^ message[348] ^ message[351] ^ message[354] ^ message[358] ^ message[361] ^ message[363] ^ message[364] ^ message[366] ^ message[367] ^ message[370] ^ message[372] ^ message[373] ^ message[376] ^ message[379] ^ message[382] ^ message[383] ^ message[386] ^ message[389] ^ message[393] ^ message[397] ^ message[398] ^ message[401] ^ message[404] ^ message[408] ^ message[413] ^ message[417] ^ message[418] ^ message[420] ^ message[421] ^ message[422] ^ message[424] ^ message[425] ^ message[427] ^ message[428] ^ message[431] ^ message[432] ^ message[434] ^ message[435] ^ message[437] ^ message[438] ^ message[441] ^ message[443] ^ message[444] ^ message[447] ^ message[450] ^ message[452] ^ message[454] ^ message[455] ^ message[457] ^ message[458] ^ message[461] ^ message[463] ^ message[464] ^ message[467] ^ message[470] ^ message[473] ^ message[474] ^ message[477] ^ message[480] ^ message[484] ^ message[487] ^ message[489] ^ message[490] ^ message[492] ^ message[493] ^ message[496] ^ message[498] ^ message[499] ^ message[502] ^ message[505] ^ message[508] ^ message[509];
    assign parity[9] = message[0] ^ message[1] ^ message[3] ^ message[4] ^ message[6] ^ message[8] ^ message[10] ^ message[12] ^ message[14] ^ message[17] ^ message[20] ^ message[22] ^ message[24] ^ message[27] ^ message[31] ^ message[35] ^ message[37] ^ message[39] ^ message[42] ^ message[46] ^ message[51] ^ message[56] ^ message[58] ^ message[60] ^ message[63] ^ message[67] ^ message[72] ^ message[78] ^ message[84] ^ message[86] ^ message[88] ^ message[91] ^ message[95] ^ message[100] ^ message[106] ^ message[113] ^ message[120] ^ message[122] ^ message[124] ^ message[127] ^ message[131] ^ message[136] ^ message[142] ^ message[149] ^ message[157] ^ message[165] ^ message[166] ^ message[167] ^ message[168] ^ message[170] ^ message[171] ^ message[172] ^ message[173] ^ message[175] ^ message[176] ^ message[177] ^ message[179] ^ message[180] ^ message[182] ^ message[184] ^ message[186] ^ message[187] ^ message[188] ^ message[190] ^ message[191] ^ message[192] ^ message[194] ^ message[195] ^ message[197] ^ message[199] ^ message[201] ^ message[202] ^ message[204] ^ message[205] ^ message[207] ^ message[209] ^ message[211] ^ message[213] ^ message[215] ^ message[218] ^ message[221] ^ message[222] ^ message[223] ^ message[225] ^ message[226] ^ message[227] ^ message[229] ^ message[230] ^ message[232] ^ message[234] ^ message[236] ^ message[237] ^ message[239] ^ message[240] ^ message[242] ^ message[244] ^ message[246] ^ message[248] ^ message[250] ^ message[253] ^ message[256] ^ message[257] ^ message[259] ^ message[260] ^ message[262] ^ message[264] ^ message[266] ^ message[268] ^ message[270] ^ message[273] ^ message[276] ^ message[278] ^ message[280] ^ message[283] ^ message[287] ^ message[291] ^ message[292] ^ message[293] ^ message[295] ^ message[296] ^ message[297] ^ message[299] ^ message[300] ^ message[302] ^ message[304] ^ message[306] ^ message[307] ^ message[309] ^ message[310] ^ message[312] ^ message[314] ^ message[316] ^ message[318] ^ message[320] ^ message[323] ^ message[326] ^ message[327] ^ message[329] ^ message[330] ^ message[332] ^ message[334] ^ message[336] ^ message[338] ^ message[340] ^ message[343] ^ message[346] ^ message[348] ^ message[350] ^ message[353] ^ message[357] ^ message[361] ^ message[362] ^ message[364] ^ message[365] ^ message[367] ^ message[369] ^ message[371] ^ message[373] ^ message[375] ^ message[378] ^ message[381] ^ message[383] ^ message[385] ^ message[388] ^ message[392] ^ message[396] ^ message[398] ^ message[400] ^ message[403] ^ message[407] ^ message[412] ^ message[417] ^ message[418] ^ message[419] ^ message[421] ^ message[422] ^ message[423] ^ message[425] ^ message[426] ^ message[428] ^ message[430] ^ message[432] ^ message[433] ^ message[435] ^ message[436] ^ message[438] ^ message[440] ^ message[442] ^ message[444] ^ message[446] ^ message[449] ^ message[452] ^ message[453] ^ message[455] ^ message[456] ^ message[458] ^ message[460] ^ message[462] ^ message[464] ^ message[466] ^ message[469] ^ message[472] ^ message[474] ^ message[476] ^ message[479] ^ message[483] ^ message[487] ^ message[488] ^ message[490] ^ message[491] ^ message[493] ^ message[495] ^ message[497] ^ message[499] ^ message[501] ^ message[504] ^ message[507] ^ message[509] ^ message[511];
    assign parity[10] = message[0] ^ message[1] ^ message[2] ^ message[4] ^ message[5] ^ message[7] ^ message[10] ^ message[11] ^ message[13] ^ message[16] ^ message[20] ^ message[21] ^ message[23] ^ message[26] ^ message[30] ^ message[35] ^ message[36] ^ message[38] ^ message[41] ^ message[45] ^ message[50] ^ message[56] ^ message[57] ^ message[59] ^ message[62] ^ message[66] ^ message[71] ^ message[77] ^ message[84] ^ message[85] ^ message[87] ^ message[90] ^ message[94] ^ message[99] ^ message[105] ^ message[112] ^ message[120] ^ message[121] ^ message[123] ^ message[126] ^ message[130] ^ message[135] ^ message[141] ^ message[148] ^ message[156] ^ message[165] ^ message[166] ^ message[167] ^ message[168] ^ message[169] ^ message[171] ^ message[172] ^ message[173] ^ message[174] ^ message[176] ^ message[177] ^ message[178] ^ message[180] ^ message[181] ^ message[183] ^ message[186] ^ message[187] ^ message[188] ^ message[189] ^ message[191] ^ message[192] ^ message[193] ^ message[195] ^ message[196] ^ message[198] ^ message[201] ^ message[202] ^ message[203] ^ message[205] ^ message[206] ^ message[208] ^ message[211] ^ message[212] ^ message[214] ^ message[217] ^ message[221] ^ message[222] ^ message[223] ^ message[224] ^ message[226] ^ message[227] ^ message[228] ^ message[230] ^ message[231] ^ message[233] ^ message[236] ^ message[237] ^ message[238] ^ message[240] ^ message[241] ^ message[243] ^ message[246] ^ message[247] ^ message[249] ^ message[252] ^ message[256] ^ message[257] ^ message[258] ^ message[260] ^ message[261] ^ message[263] ^ message[266] ^ message[267] ^ message[269] ^ message[272] ^ message[276] ^ message[277] ^ message[279] ^ message[282] ^ message[286] ^ message[291] ^ message[292] ^ message[293] ^ message[294] ^ message[296] ^ message[297] ^ message[298] ^ message[300] ^ message[301] ^ message[303] ^ message[306] ^ message[307] ^ message[308] ^ message[310] ^ message[311] ^ message[313] ^ message[316] ^ message[317] ^ message[319] ^ message[322] ^ message[326] ^ message[327] ^ message[328] ^ message[330] ^ message[331] ^ message[333] ^ message[336] ^ message[337] ^ message[339] ^ message[342] ^ message[346] ^ message[347] ^ message[349] ^ message[352] ^ message[356] ^ message[361] ^ message[362] ^ message[363] ^ message[365] ^ message[366] ^ message[368] ^ message[371] ^ message[372] ^ message[374] ^ message[377] ^ message[381] ^ message[382] ^ message[384] ^ message[387] ^ message[391] ^ message[396] ^ message[397] ^ message[399] ^ message[402] ^ message[406] ^ message[411] ^ message[417] ^ message[418] ^ message[419] ^ message[420] ^ message[422] ^ message[423] ^ message[424] ^ message[426] ^ message[427] ^ message[429] ^ message[432] ^ message[433] ^ message[434] ^ message[436] ^ message[437] ^ message[439] ^ message[442] ^ message[443] ^ message[445] ^ message[448] ^ message[452] ^ message[453] ^ message[454] ^ message[456] ^ message[457] ^ message[459] ^ message[462] ^ message[463] ^ message[465] ^ message[468] ^ message[472] ^ message[473] ^ message[475] ^ message[478] ^ message[482] ^ message[487] ^ message[488] ^ message[489] ^ message[491] ^ message[492] ^ message[494] ^ message[497] ^ message[498] ^ message[500] ^ message[503] ^ message[507] ^ message[508] ^ message[510];
  end else if ((CodewordWidth == 1036) && (MessageWidth == 1024)) begin : gen_1036_1024
    `BR_ASSERT_STATIC(parity_width_matches_a, ParityWidth == 12)
    assign parity[0] = message[165] ^ message[166] ^ message[167] ^ message[168] ^ message[169] ^ message[170] ^ message[171] ^ message[172] ^ message[173] ^ message[174] ^ message[175] ^ message[176] ^ message[177] ^ message[178] ^ message[179] ^ message[180] ^ message[181] ^ message[182] ^ message[183] ^ message[184] ^ message[185] ^ message[186] ^ message[187] ^ message[188] ^ message[189] ^ message[190] ^ message[191] ^ message[192] ^ message[193] ^ message[194] ^ message[195] ^ message[196] ^ message[197] ^ message[198] ^ message[199] ^ message[200] ^ message[201] ^ message[202] ^ message[203] ^ message[204] ^ message[205] ^ message[206] ^ message[207] ^ message[208] ^ message[209] ^ message[210] ^ message[211] ^ message[212] ^ message[213] ^ message[214] ^ message[215] ^ message[216] ^ message[217] ^ message[218] ^ message[219] ^ message[682] ^ message[683] ^ message[684] ^ message[685] ^ message[686] ^ message[687] ^ message[688] ^ message[689] ^ message[690] ^ message[691] ^ message[692] ^ message[693] ^ message[694] ^ message[695] ^ message[696] ^ message[697] ^ message[698] ^ message[699] ^ message[700] ^ message[701] ^ message[702] ^ message[703] ^ message[704] ^ message[705] ^ message[706] ^ message[707] ^ message[708] ^ message[709] ^ message[710] ^ message[711] ^ message[712] ^ message[713] ^ message[714] ^ message[715] ^ message[716] ^ message[717] ^ message[718] ^ message[719] ^ message[720] ^ message[721] ^ message[722] ^ message[723] ^ message[724] ^ message[725] ^ message[726] ^ message[727] ^ message[728] ^ message[729] ^ message[730] ^ message[731] ^ message[732] ^ message[733] ^ message[734] ^ message[735] ^ message[736] ^ message[737] ^ message[738] ^ message[739] ^ message[740] ^ message[741] ^ message[742] ^ message[743] ^ message[744] ^ message[745] ^ message[746] ^ message[747] ^ message[748] ^ message[749] ^ message[750] ^ message[751] ^ message[752] ^ message[753] ^ message[754] ^ message[755] ^ message[756] ^ message[757] ^ message[758] ^ message[759] ^ message[760] ^ message[761] ^ message[762] ^ message[763] ^ message[764] ^ message[765] ^ message[766] ^ message[767] ^ message[768] ^ message[769] ^ message[770] ^ message[771] ^ message[772] ^ message[773] ^ message[774] ^ message[775] ^ message[776] ^ message[777] ^ message[778] ^ message[779] ^ message[780] ^ message[781] ^ message[782] ^ message[783] ^ message[784] ^ message[785] ^ message[786] ^ message[787] ^ message[788] ^ message[789] ^ message[790] ^ message[791] ^ message[792] ^ message[793] ^ message[794] ^ message[795] ^ message[796] ^ message[797] ^ message[798] ^ message[799] ^ message[800] ^ message[801] ^ message[802] ^ message[803] ^ message[804] ^ message[805] ^ message[806] ^ message[807] ^ message[808] ^ message[809] ^ message[810] ^ message[811] ^ message[812] ^ message[813] ^ message[814] ^ message[815] ^ message[816] ^ message[817] ^ message[818] ^ message[819] ^ message[820] ^ message[821] ^ message[822] ^ message[823] ^ message[824] ^ message[825] ^ message[826] ^ message[827] ^ message[828] ^ message[829] ^ message[830] ^ message[831] ^ message[832] ^ message[833] ^ message[834] ^ message[835] ^ message[836] ^ message[837] ^ message[838] ^ message[839] ^ message[840] ^ message[841] ^ message[842] ^ message[843] ^ message[844] ^ message[845] ^ message[846] ^ message[847] ^ message[848] ^ message[849] ^ message[850] ^ message[851] ^ message[852] ^ message[853] ^ message[854] ^ message[855] ^ message[856] ^ message[857] ^ message[858] ^ message[859] ^ message[860] ^ message[861] ^ message[862] ^ message[863] ^ message[864] ^ message[865] ^ message[866] ^ message[867] ^ message[868] ^ message[869] ^ message[870] ^ message[871] ^ message[872] ^ message[873] ^ message[874] ^ message[875] ^ message[876] ^ message[877] ^ message[878] ^ message[879] ^ message[880] ^ message[881] ^ message[882] ^ message[883] ^ message[884] ^ message[885] ^ message[886] ^ message[887] ^ message[888] ^ message[889] ^ message[890] ^ message[891] ^ message[892] ^ message[893] ^ message[894] ^ message[895] ^ message[896] ^ message[897] ^ message[898] ^ message[899] ^ message[900] ^ message[901] ^ message[902] ^ message[903] ^ message[904] ^ message[905] ^ message[906] ^ message[907] ^ message[908] ^ message[909] ^ message[910] ^ message[911] ^ message[912] ^ message[913] ^ message[914] ^ message[915] ^ message[916] ^ message[917] ^ message[918] ^ message[919] ^ message[920] ^ message[921] ^ message[922] ^ message[923] ^ message[924] ^ message[925] ^ message[926] ^ message[927] ^ message[928] ^ message[929] ^ message[930] ^ message[931] ^ message[932] ^ message[933] ^ message[934] ^ message[935] ^ message[936] ^ message[937] ^ message[938] ^ message[939] ^ message[940] ^ message[941] ^ message[942] ^ message[943] ^ message[944] ^ message[945] ^ message[946] ^ message[947] ^ message[948] ^ message[949] ^ message[950] ^ message[951] ^ message[952] ^ message[953] ^ message[954] ^ message[955] ^ message[956] ^ message[957] ^ message[958] ^ message[959] ^ message[960] ^ message[961] ^ message[962] ^ message[963] ^ message[964] ^ message[965] ^ message[966] ^ message[967] ^ message[968] ^ message[969] ^ message[970] ^ message[971] ^ message[972] ^ message[973] ^ message[974] ^ message[975] ^ message[976] ^ message[977] ^ message[978] ^ message[979] ^ message[980] ^ message[981] ^ message[982] ^ message[983] ^ message[984] ^ message[985] ^ message[986] ^ message[987] ^ message[988] ^ message[989] ^ message[990] ^ message[991] ^ message[992] ^ message[993] ^ message[994] ^ message[995] ^ message[996] ^ message[997] ^ message[998] ^ message[999] ^ message[1000] ^ message[1001] ^ message[1002] ^ message[1003] ^ message[1004] ^ message[1005] ^ message[1006] ^ message[1007] ^ message[1008] ^ message[1009] ^ message[1010] ^ message[1011];
    assign parity[1] = message[120] ^ message[121] ^ message[122] ^ message[123] ^ message[124] ^ message[125] ^ message[126] ^ message[127] ^ message[128] ^ message[129] ^ message[130] ^ message[131] ^ message[132] ^ message[133] ^ message[134] ^ message[135] ^ message[136] ^ message[137] ^ message[138] ^ message[139] ^ message[140] ^ message[141] ^ message[142] ^ message[143] ^ message[144] ^ message[145] ^ message[146] ^ message[147] ^ message[148] ^ message[149] ^ message[150] ^ message[151] ^ message[152] ^ message[153] ^ message[154] ^ message[155] ^ message[156] ^ message[157] ^ message[158] ^ message[159] ^ message[160] ^ message[161] ^ message[162] ^ message[163] ^ message[164] ^ message[210] ^ message[211] ^ message[212] ^ message[213] ^ message[214] ^ message[215] ^ message[216] ^ message[217] ^ message[218] ^ message[219] ^ message[472] ^ message[473] ^ message[474] ^ message[475] ^ message[476] ^ message[477] ^ message[478] ^ message[479] ^ message[480] ^ message[481] ^ message[482] ^ message[483] ^ message[484] ^ message[485] ^ message[486] ^ message[487] ^ message[488] ^ message[489] ^ message[490] ^ message[491] ^ message[492] ^ message[493] ^ message[494] ^ message[495] ^ message[496] ^ message[497] ^ message[498] ^ message[499] ^ message[500] ^ message[501] ^ message[502] ^ message[503] ^ message[504] ^ message[505] ^ message[506] ^ message[507] ^ message[508] ^ message[509] ^ message[510] ^ message[511] ^ message[512] ^ message[513] ^ message[514] ^ message[515] ^ message[516] ^ message[517] ^ message[518] ^ message[519] ^ message[520] ^ message[521] ^ message[522] ^ message[523] ^ message[524] ^ message[525] ^ message[526] ^ message[527] ^ message[528] ^ message[529] ^ message[530] ^ message[531] ^ message[532] ^ message[533] ^ message[534] ^ message[535] ^ message[536] ^ message[537] ^ message[538] ^ message[539] ^ message[540] ^ message[541] ^ message[542] ^ message[543] ^ message[544] ^ message[545] ^ message[546] ^ message[547] ^ message[548] ^ message[549] ^ message[550] ^ message[551] ^ message[552] ^ message[553] ^ message[554] ^ message[555] ^ message[556] ^ message[557] ^ message[558] ^ message[559] ^ message[560] ^ message[561] ^ message[562] ^ message[563] ^ message[564] ^ message[565] ^ message[566] ^ message[567] ^ message[568] ^ message[569] ^ message[570] ^ message[571] ^ message[572] ^ message[573] ^ message[574] ^ message[575] ^ message[576] ^ message[577] ^ message[578] ^ message[579] ^ message[580] ^ message[581] ^ message[582] ^ message[583] ^ message[584] ^ message[585] ^ message[586] ^ message[587] ^ message[588] ^ message[589] ^ message[590] ^ message[591] ^ message[592] ^ message[593] ^ message[594] ^ message[595] ^ message[596] ^ message[597] ^ message[598] ^ message[599] ^ message[600] ^ message[601] ^ message[602] ^ message[603] ^ message[604] ^ message[605] ^ message[606] ^ message[607] ^ message[608] ^ message[609] ^ message[610] ^ message[611] ^ message[612] ^ message[613] ^ message[614] ^ message[615] ^ message[616] ^ message[617] ^ message[618] ^ message[619] ^ message[620] ^ message[621] ^ message[622] ^ message[623] ^ message[624] ^ message[625] ^ message[626] ^ message[627] ^ message[628] ^ message[629] ^ message[630] ^ message[631] ^ message[632] ^ message[633] ^ message[634] ^ message[635] ^ message[636] ^ message[637] ^ message[638] ^ message[639] ^ message[640] ^ message[641] ^ message[642] ^ message[643] ^ message[644] ^ message[645] ^ message[646] ^ message[647] ^ message[648] ^ message[649] ^ message[650] ^ message[651] ^ message[652] ^ message[653] ^ message[654] ^ message[655] ^ message[656] ^ message[657] ^ message[658] ^ message[659] ^ message[660] ^ message[661] ^ message[662] ^ message[663] ^ message[664] ^ message[665] ^ message[666] ^ message[667] ^ message[668] ^ message[669] ^ message[670] ^ message[671] ^ message[672] ^ message[673] ^ message[674] ^ message[675] ^ message[676] ^ message[677] ^ message[678] ^ message[679] ^ message[680] ^ message[681] ^ message[892] ^ message[893] ^ message[894] ^ message[895] ^ message[896] ^ message[897] ^ message[898] ^ message[899] ^ message[900] ^ message[901] ^ message[902] ^ message[903] ^ message[904] ^ message[905] ^ message[906] ^ message[907] ^ message[908] ^ message[909] ^ message[910] ^ message[911] ^ message[912] ^ message[913] ^ message[914] ^ message[915] ^ message[916] ^ message[917] ^ message[918] ^ message[919] ^ message[920] ^ message[921] ^ message[922] ^ message[923] ^ message[924] ^ message[925] ^ message[926] ^ message[927] ^ message[928] ^ message[929] ^ message[930] ^ message[931] ^ message[932] ^ message[933] ^ message[934] ^ message[935] ^ message[936] ^ message[937] ^ message[938] ^ message[939] ^ message[940] ^ message[941] ^ message[942] ^ message[943] ^ message[944] ^ message[945] ^ message[946] ^ message[947] ^ message[948] ^ message[949] ^ message[950] ^ message[951] ^ message[952] ^ message[953] ^ message[954] ^ message[955] ^ message[956] ^ message[957] ^ message[958] ^ message[959] ^ message[960] ^ message[961] ^ message[962] ^ message[963] ^ message[964] ^ message[965] ^ message[966] ^ message[967] ^ message[968] ^ message[969] ^ message[970] ^ message[971] ^ message[972] ^ message[973] ^ message[974] ^ message[975] ^ message[976] ^ message[977] ^ message[978] ^ message[979] ^ message[980] ^ message[981] ^ message[982] ^ message[983] ^ message[984] ^ message[985] ^ message[986] ^ message[987] ^ message[988] ^ message[989] ^ message[990] ^ message[991] ^ message[992] ^ message[993] ^ message[994] ^ message[995] ^ message[996] ^ message[997] ^ message[998] ^ message[999] ^ message[1000] ^ message[1001] ^ message[1002] ^ message[1003] ^ message[1004] ^ message[1005] ^ message[1006] ^ message[1007] ^ message[1008] ^ message[1009] ^ message[1010] ^ message[1011];
    assign parity[2] = message[84] ^ message[85] ^ message[86] ^ message[87] ^ message[88] ^ message[89] ^ message[90] ^ message[91] ^ message[92] ^ message[93] ^ message[94] ^ message[95] ^ message[96] ^ message[97] ^ message[98] ^ message[99] ^ message[100] ^ message[101] ^ message[102] ^ message[103] ^ message[104] ^ message[105] ^ message[106] ^ message[107] ^ message[108] ^ message[109] ^ message[110] ^ message[111] ^ message[112] ^ message[113] ^ message[114] ^ message[115] ^ message[116] ^ message[117] ^ message[118] ^ message[119] ^ message[156] ^ message[157] ^ message[158] ^ message[159] ^ message[160] ^ message[161] ^ message[162] ^ message[163] ^ message[164] ^ message[201] ^ message[202] ^ message[203] ^ message[204] ^ message[205] ^ message[206] ^ message[207] ^ message[208] ^ message[209] ^ message[219] ^ message[346] ^ message[347] ^ message[348] ^ message[349] ^ message[350] ^ message[351] ^ message[352] ^ message[353] ^ message[354] ^ message[355] ^ message[356] ^ message[357] ^ message[358] ^ message[359] ^ message[360] ^ message[361] ^ message[362] ^ message[363] ^ message[364] ^ message[365] ^ message[366] ^ message[367] ^ message[368] ^ message[369] ^ message[370] ^ message[371] ^ message[372] ^ message[373] ^ message[374] ^ message[375] ^ message[376] ^ message[377] ^ message[378] ^ message[379] ^ message[380] ^ message[381] ^ message[382] ^ message[383] ^ message[384] ^ message[385] ^ message[386] ^ message[387] ^ message[388] ^ message[389] ^ message[390] ^ message[391] ^ message[392] ^ message[393] ^ message[394] ^ message[395] ^ message[396] ^ message[397] ^ message[398] ^ message[399] ^ message[400] ^ message[401] ^ message[402] ^ message[403] ^ message[404] ^ message[405] ^ message[406] ^ message[407] ^ message[408] ^ message[409] ^ message[410] ^ message[411] ^ message[412] ^ message[413] ^ message[414] ^ message[415] ^ message[416] ^ message[417] ^ message[418] ^ message[419] ^ message[420] ^ message[421] ^ message[422] ^ message[423] ^ message[424] ^ message[425] ^ message[426] ^ message[427] ^ message[428] ^ message[429] ^ message[430] ^ message[431] ^ message[432] ^ message[433] ^ message[434] ^ message[435] ^ message[436] ^ message[437] ^ message[438] ^ message[439] ^ message[440] ^ message[441] ^ message[442] ^ message[443] ^ message[444] ^ message[445] ^ message[446] ^ message[447] ^ message[448] ^ message[449] ^ message[450] ^ message[451] ^ message[452] ^ message[453] ^ message[454] ^ message[455] ^ message[456] ^ message[457] ^ message[458] ^ message[459] ^ message[460] ^ message[461] ^ message[462] ^ message[463] ^ message[464] ^ message[465] ^ message[466] ^ message[467] ^ message[468] ^ message[469] ^ message[470] ^ message[471] ^ message[598] ^ message[599] ^ message[600] ^ message[601] ^ message[602] ^ message[603] ^ message[604] ^ message[605] ^ message[606] ^ message[607] ^ message[608] ^ message[609] ^ message[610] ^ message[611] ^ message[612] ^ message[613] ^ message[614] ^ message[615] ^ message[616] ^ message[617] ^ message[618] ^ message[619] ^ message[620] ^ message[621] ^ message[622] ^ message[623] ^ message[624] ^ message[625] ^ message[626] ^ message[627] ^ message[628] ^ message[629] ^ message[630] ^ message[631] ^ message[632] ^ message[633] ^ message[634] ^ message[635] ^ message[636] ^ message[637] ^ message[638] ^ message[639] ^ message[640] ^ message[641] ^ message[642] ^ message[643] ^ message[644] ^ message[645] ^ message[646] ^ message[647] ^ message[648] ^ message[649] ^ message[650] ^ message[651] ^ message[652] ^ message[653] ^ message[654] ^ message[655] ^ message[656] ^ message[657] ^ message[658] ^ message[659] ^ message[660] ^ message[661] ^ message[662] ^ message[663] ^ message[664] ^ message[665] ^ message[666] ^ message[667] ^ message[668] ^ message[669] ^ message[670] ^ message[671] ^ message[672] ^ message[673] ^ message[674] ^ message[675] ^ message[676] ^ message[677] ^ message[678] ^ message[679] ^ message[680] ^ message[681] ^ message[808] ^ message[809] ^ message[810] ^ message[811] ^ message[812] ^ message[813] ^ message[814] ^ message[815] ^ message[816] ^ message[817] ^ message[818] ^ message[819] ^ message[820] ^ message[821] ^ message[822] ^ message[823] ^ message[824] ^ message[825] ^ message[826] ^ message[827] ^ message[828] ^ message[829] ^ message[830] ^ message[831] ^ message[832] ^ message[833] ^ message[834] ^ message[835] ^ message[836] ^ message[837] ^ message[838] ^ message[839] ^ message[840] ^ message[841] ^ message[842] ^ message[843] ^ message[844] ^ message[845] ^ message[846] ^ message[847] ^ message[848] ^ message[849] ^ message[850] ^ message[851] ^ message[852] ^ message[853] ^ message[854] ^ message[855] ^ message[856] ^ message[857] ^ message[858] ^ message[859] ^ message[860] ^ message[861] ^ message[862] ^ message[863] ^ message[864] ^ message[865] ^ message[866] ^ message[867] ^ message[868] ^ message[869] ^ message[870] ^ message[871] ^ message[872] ^ message[873] ^ message[874] ^ message[875] ^ message[876] ^ message[877] ^ message[878] ^ message[879] ^ message[880] ^ message[881] ^ message[882] ^ message[883] ^ message[884] ^ message[885] ^ message[886] ^ message[887] ^ message[888] ^ message[889] ^ message[890] ^ message[891] ^ message[976] ^ message[977] ^ message[978] ^ message[979] ^ message[980] ^ message[981] ^ message[982] ^ message[983] ^ message[984] ^ message[985] ^ message[986] ^ message[987] ^ message[988] ^ message[989] ^ message[990] ^ message[991] ^ message[992] ^ message[993] ^ message[994] ^ message[995] ^ message[996] ^ message[997] ^ message[998] ^ message[999] ^ message[1000] ^ message[1001] ^ message[1002] ^ message[1003] ^ message[1004] ^ message[1005] ^ message[1006] ^ message[1007] ^ message[1008] ^ message[1009] ^ message[1010] ^ message[1011];
    assign parity[3] = message[56] ^ message[57] ^ message[58] ^ message[59] ^ message[60] ^ message[61] ^ message[62] ^ message[63] ^ message[64] ^ message[65] ^ message[66] ^ message[67] ^ message[68] ^ message[69] ^ message[70] ^ message[71] ^ message[72] ^ message[73] ^ message[74] ^ message[75] ^ message[76] ^ message[77] ^ message[78] ^ message[79] ^ message[80] ^ message[81] ^ message[82] ^ message[83] ^ message[112] ^ message[113] ^ message[114] ^ message[115] ^ message[116] ^ message[117] ^ message[118] ^ message[119] ^ message[148] ^ message[149] ^ message[150] ^ message[151] ^ message[152] ^ message[153] ^ message[154] ^ message[155] ^ message[164] ^ message[193] ^ message[194] ^ message[195] ^ message[196] ^ message[197] ^ message[198] ^ message[199] ^ message[200] ^ message[209] ^ message[218] ^ message[276] ^ message[277] ^ message[278] ^ message[279] ^ message[280] ^ message[281] ^ message[282] ^ message[283] ^ message[284] ^ message[285] ^ message[286] ^ message[287] ^ message[288] ^ message[289] ^ message[290] ^ message[291] ^ message[292] ^ message[293] ^ message[294] ^ message[295] ^ message[296] ^ message[297] ^ message[298] ^ message[299] ^ message[300] ^ message[301] ^ message[302] ^ message[303] ^ message[304] ^ message[305] ^ message[306] ^ message[307] ^ message[308] ^ message[309] ^ message[310] ^ message[311] ^ message[312] ^ message[313] ^ message[314] ^ message[315] ^ message[316] ^ message[317] ^ message[318] ^ message[319] ^ message[320] ^ message[321] ^ message[322] ^ message[323] ^ message[324] ^ message[325] ^ message[326] ^ message[327] ^ message[328] ^ message[329] ^ message[330] ^ message[331] ^ message[332] ^ message[333] ^ message[334] ^ message[335] ^ message[336] ^ message[337] ^ message[338] ^ message[339] ^ message[340] ^ message[341] ^ message[342] ^ message[343] ^ message[344] ^ message[345] ^ message[416] ^ message[417] ^ message[418] ^ message[419] ^ message[420] ^ message[421] ^ message[422] ^ message[423] ^ message[424] ^ message[425] ^ message[426] ^ message[427] ^ message[428] ^ message[429] ^ message[430] ^ message[431] ^ message[432] ^ message[433] ^ message[434] ^ message[435] ^ message[436] ^ message[437] ^ message[438] ^ message[439] ^ message[440] ^ message[441] ^ message[442] ^ message[443] ^ message[444] ^ message[445] ^ message[446] ^ message[447] ^ message[448] ^ message[449] ^ message[450] ^ message[451] ^ message[452] ^ message[453] ^ message[454] ^ message[455] ^ message[456] ^ message[457] ^ message[458] ^ message[459] ^ message[460] ^ message[461] ^ message[462] ^ message[463] ^ message[464] ^ message[465] ^ message[466] ^ message[467] ^ message[468] ^ message[469] ^ message[470] ^ message[471] ^ message[542] ^ message[543] ^ message[544] ^ message[545] ^ message[546] ^ message[547] ^ message[548] ^ message[549] ^ message[550] ^ message[551] ^ message[552] ^ message[553] ^ message[554] ^ message[555] ^ message[556] ^ message[557] ^ message[558] ^ message[559] ^ message[560] ^ message[561] ^ message[562] ^ message[563] ^ message[564] ^ message[565] ^ message[566] ^ message[567] ^ message[568] ^ message[569] ^ message[570] ^ message[571] ^ message[572] ^ message[573] ^ message[574] ^ message[575] ^ message[576] ^ message[577] ^ message[578] ^ message[579] ^ message[580] ^ message[581] ^ message[582] ^ message[583] ^ message[584] ^ message[585] ^ message[586] ^ message[587] ^ message[588] ^ message[589] ^ message[590] ^ message[591] ^ message[592] ^ message[593] ^ message[594] ^ message[595] ^ message[596] ^ message[597] ^ message[654] ^ message[655] ^ message[656] ^ message[657] ^ message[658] ^ message[659] ^ message[660] ^ message[661] ^ message[662] ^ message[663] ^ message[664] ^ message[665] ^ message[666] ^ message[667] ^ message[668] ^ message[669] ^ message[670] ^ message[671] ^ message[672] ^ message[673] ^ message[674] ^ message[675] ^ message[676] ^ message[677] ^ message[678] ^ message[679] ^ message[680] ^ message[681] ^ message[752] ^ message[753] ^ message[754] ^ message[755] ^ message[756] ^ message[757] ^ message[758] ^ message[759] ^ message[760] ^ message[761] ^ message[762] ^ message[763] ^ message[764] ^ message[765] ^ message[766] ^ message[767] ^ message[768] ^ message[769] ^ message[770] ^ message[771] ^ message[772] ^ message[773] ^ message[774] ^ message[775] ^ message[776] ^ message[777] ^ message[778] ^ message[779] ^ message[780] ^ message[781] ^ message[782] ^ message[783] ^ message[784] ^ message[785] ^ message[786] ^ message[787] ^ message[788] ^ message[789] ^ message[790] ^ message[791] ^ message[792] ^ message[793] ^ message[794] ^ message[795] ^ message[796] ^ message[797] ^ message[798] ^ message[799] ^ message[800] ^ message[801] ^ message[802] ^ message[803] ^ message[804] ^ message[805] ^ message[806] ^ message[807] ^ message[864] ^ message[865] ^ message[866] ^ message[867] ^ message[868] ^ message[869] ^ message[870] ^ message[871] ^ message[872] ^ message[873] ^ message[874] ^ message[875] ^ message[876] ^ message[877] ^ message[878] ^ message[879] ^ message[880] ^ message[881] ^ message[882] ^ message[883] ^ message[884] ^ message[885] ^ message[886] ^ message[887] ^ message[888] ^ message[889] ^ message[890] ^ message[891] ^ message[948] ^ message[949] ^ message[950] ^ message[951] ^ message[952] ^ message[953] ^ message[954] ^ message[955] ^ message[956] ^ message[957] ^ message[958] ^ message[959] ^ message[960] ^ message[961] ^ message[962] ^ message[963] ^ message[964] ^ message[965] ^ message[966] ^ message[967] ^ message[968] ^ message[969] ^ message[970] ^ message[971] ^ message[972] ^ message[973] ^ message[974] ^ message[975] ^ message[1004] ^ message[1005] ^ message[1006] ^ message[1007] ^ message[1008] ^ message[1009] ^ message[1010] ^ message[1011] ^ message[1020] ^ message[1021] ^ message[1022] ^ message[1023];
    assign parity[4] = message[35] ^ message[36] ^ message[37] ^ message[38] ^ message[39] ^ message[40] ^ message[41] ^ message[42] ^ message[43] ^ message[44] ^ message[45] ^ message[46] ^ message[47] ^ message[48] ^ message[49] ^ message[50] ^ message[51] ^ message[52] ^ message[53] ^ message[54] ^ message[55] ^ message[77] ^ message[78] ^ message[79] ^ message[80] ^ message[81] ^ message[82] ^ message[83] ^ message[105] ^ message[106] ^ message[107] ^ message[108] ^ message[109] ^ message[110] ^ message[111] ^ message[119] ^ message[141] ^ message[142] ^ message[143] ^ message[144] ^ message[145] ^ message[146] ^ message[147] ^ message[155] ^ message[163] ^ message[186] ^ message[187] ^ message[188] ^ message[189] ^ message[190] ^ message[191] ^ message[192] ^ message[200] ^ message[208] ^ message[217] ^ message[241] ^ message[242] ^ message[243] ^ message[244] ^ message[245] ^ message[246] ^ message[247] ^ message[248] ^ message[249] ^ message[250] ^ message[251] ^ message[252] ^ message[253] ^ message[254] ^ message[255] ^ message[256] ^ message[257] ^ message[258] ^ message[259] ^ message[260] ^ message[261] ^ message[262] ^ message[263] ^ message[264] ^ message[265] ^ message[266] ^ message[267] ^ message[268] ^ message[269] ^ message[270] ^ message[271] ^ message[272] ^ message[273] ^ message[274] ^ message[275] ^ message[311] ^ message[312] ^ message[313] ^ message[314] ^ message[315] ^ message[316] ^ message[317] ^ message[318] ^ message[319] ^ message[320] ^ message[321] ^ message[322] ^ message[323] ^ message[324] ^ message[325] ^ message[326] ^ message[327] ^ message[328] ^ message[329] ^ message[330] ^ message[331] ^ message[332] ^ message[333] ^ message[334] ^ message[335] ^ message[336] ^ message[337] ^ message[338] ^ message[339] ^ message[340] ^ message[341] ^ message[342] ^ message[343] ^ message[344] ^ message[345] ^ message[381] ^ message[382] ^ message[383] ^ message[384] ^ message[385] ^ message[386] ^ message[387] ^ message[388] ^ message[389] ^ message[390] ^ message[391] ^ message[392] ^ message[393] ^ message[394] ^ message[395] ^ message[396] ^ message[397] ^ message[398] ^ message[399] ^ message[400] ^ message[401] ^ message[402] ^ message[403] ^ message[404] ^ message[405] ^ message[406] ^ message[407] ^ message[408] ^ message[409] ^ message[410] ^ message[411] ^ message[412] ^ message[413] ^ message[414] ^ message[415] ^ message[451] ^ message[452] ^ message[453] ^ message[454] ^ message[455] ^ message[456] ^ message[457] ^ message[458] ^ message[459] ^ message[460] ^ message[461] ^ message[462] ^ message[463] ^ message[464] ^ message[465] ^ message[466] ^ message[467] ^ message[468] ^ message[469] ^ message[470] ^ message[471] ^ message[507] ^ message[508] ^ message[509] ^ message[510] ^ message[511] ^ message[512] ^ message[513] ^ message[514] ^ message[515] ^ message[516] ^ message[517] ^ message[518] ^ message[519] ^ message[520] ^ message[521] ^ message[522] ^ message[523] ^ message[524] ^ message[525] ^ message[526] ^ message[527] ^ message[528] ^ message[529] ^ message[530] ^ message[531] ^ message[532] ^ message[533] ^ message[534] ^ message[535] ^ message[536] ^ message[537] ^ message[538] ^ message[539] ^ message[540] ^ message[541] ^ message[577] ^ message[578] ^ message[579] ^ message[580] ^ message[581] ^ message[582] ^ message[583] ^ message[584] ^ message[585] ^ message[586] ^ message[587] ^ message[588] ^ message[589] ^ message[590] ^ message[591] ^ message[592] ^ message[593] ^ message[594] ^ message[595] ^ message[596] ^ message[597] ^ message[633] ^ message[634] ^ message[635] ^ message[636] ^ message[637] ^ message[638] ^ message[639] ^ message[640] ^ message[641] ^ message[642] ^ message[643] ^ message[644] ^ message[645] ^ message[646] ^ message[647] ^ message[648] ^ message[649] ^ message[650] ^ message[651] ^ message[652] ^ message[653] ^ message[675] ^ message[676] ^ message[677] ^ message[678] ^ message[679] ^ message[680] ^ message[681] ^ message[717] ^ message[718] ^ message[719] ^ message[720] ^ message[721] ^ message[722] ^ message[723] ^ message[724] ^ message[725] ^ message[726] ^ message[727] ^ message[728] ^ message[729] ^ message[730] ^ message[731] ^ message[732] ^ message[733] ^ message[734] ^ message[735] ^ message[736] ^ message[737] ^ message[738] ^ message[739] ^ message[740] ^ message[741] ^ message[742] ^ message[743] ^ message[744] ^ message[745] ^ message[746] ^ message[747] ^ message[748] ^ message[749] ^ message[750] ^ message[751] ^ message[787] ^ message[788] ^ message[789] ^ message[790] ^ message[791] ^ message[792] ^ message[793] ^ message[794] ^ message[795] ^ message[796] ^ message[797] ^ message[798] ^ message[799] ^ message[800] ^ message[801] ^ message[802] ^ message[803] ^ message[804] ^ message[805] ^ message[806] ^ message[807] ^ message[843] ^ message[844] ^ message[845] ^ message[846] ^ message[847] ^ message[848] ^ message[849] ^ message[850] ^ message[851] ^ message[852] ^ message[853] ^ message[854] ^ message[855] ^ message[856] ^ message[857] ^ message[858] ^ message[859] ^ message[860] ^ message[861] ^ message[862] ^ message[863] ^ message[885] ^ message[886] ^ message[887] ^ message[888] ^ message[889] ^ message[890] ^ message[891] ^ message[927] ^ message[928] ^ message[929] ^ message[930] ^ message[931] ^ message[932] ^ message[933] ^ message[934] ^ message[935] ^ message[936] ^ message[937] ^ message[938] ^ message[939] ^ message[940] ^ message[941] ^ message[942] ^ message[943] ^ message[944] ^ message[945] ^ message[946] ^ message[947] ^ message[969] ^ message[970] ^ message[971] ^ message[972] ^ message[973] ^ message[974] ^ message[975] ^ message[997] ^ message[998] ^ message[999] ^ message[1000] ^ message[1001] ^ message[1002] ^ message[1003] ^ message[1011] ^ message[1013] ^ message[1014] ^ message[1015] ^ message[1016] ^ message[1017] ^ message[1018] ^ message[1019];
    assign parity[5] = message[20] ^ message[21] ^ message[22] ^ message[23] ^ message[24] ^ message[25] ^ message[26] ^ message[27] ^ message[28] ^ message[29] ^ message[30] ^ message[31] ^ message[32] ^ message[33] ^ message[34] ^ message[50] ^ message[51] ^ message[52] ^ message[53] ^ message[54] ^ message[55] ^ message[71] ^ message[72] ^ message[73] ^ message[74] ^ message[75] ^ message[76] ^ message[83] ^ message[99] ^ message[100] ^ message[101] ^ message[102] ^ message[103] ^ message[104] ^ message[111] ^ message[118] ^ message[135] ^ message[136] ^ message[137] ^ message[138] ^ message[139] ^ message[140] ^ message[147] ^ message[154] ^ message[162] ^ message[180] ^ message[181] ^ message[182] ^ message[183] ^ message[184] ^ message[185] ^ message[192] ^ message[199] ^ message[207] ^ message[216] ^ message[226] ^ message[227] ^ message[228] ^ message[229] ^ message[230] ^ message[231] ^ message[232] ^ message[233] ^ message[234] ^ message[235] ^ message[236] ^ message[237] ^ message[238] ^ message[239] ^ message[240] ^ message[256] ^ message[257] ^ message[258] ^ message[259] ^ message[260] ^ message[261] ^ message[262] ^ message[263] ^ message[264] ^ message[265] ^ message[266] ^ message[267] ^ message[268] ^ message[269] ^ message[270] ^ message[271] ^ message[272] ^ message[273] ^ message[274] ^ message[275] ^ message[291] ^ message[292] ^ message[293] ^ message[294] ^ message[295] ^ message[296] ^ message[297] ^ message[298] ^ message[299] ^ message[300] ^ message[301] ^ message[302] ^ message[303] ^ message[304] ^ message[305] ^ message[306] ^ message[307] ^ message[308] ^ message[309] ^ message[310] ^ message[331] ^ message[332] ^ message[333] ^ message[334] ^ message[335] ^ message[336] ^ message[337] ^ message[338] ^ message[339] ^ message[340] ^ message[341] ^ message[342] ^ message[343] ^ message[344] ^ message[345] ^ message[361] ^ message[362] ^ message[363] ^ message[364] ^ message[365] ^ message[366] ^ message[367] ^ message[368] ^ message[369] ^ message[370] ^ message[371] ^ message[372] ^ message[373] ^ message[374] ^ message[375] ^ message[376] ^ message[377] ^ message[378] ^ message[379] ^ message[380] ^ message[401] ^ message[402] ^ message[403] ^ message[404] ^ message[405] ^ message[406] ^ message[407] ^ message[408] ^ message[409] ^ message[410] ^ message[411] ^ message[412] ^ message[413] ^ message[414] ^ message[415] ^ message[436] ^ message[437] ^ message[438] ^ message[439] ^ message[440] ^ message[441] ^ message[442] ^ message[443] ^ message[444] ^ message[445] ^ message[446] ^ message[447] ^ message[448] ^ message[449] ^ message[450] ^ message[466] ^ message[467] ^ message[468] ^ message[469] ^ message[470] ^ message[471] ^ message[487] ^ message[488] ^ message[489] ^ message[490] ^ message[491] ^ message[492] ^ message[493] ^ message[494] ^ message[495] ^ message[496] ^ message[497] ^ message[498] ^ message[499] ^ message[500] ^ message[501] ^ message[502] ^ message[503] ^ message[504] ^ message[505] ^ message[506] ^ message[527] ^ message[528] ^ message[529] ^ message[530] ^ message[531] ^ message[532] ^ message[533] ^ message[534] ^ message[535] ^ message[536] ^ message[537] ^ message[538] ^ message[539] ^ message[540] ^ message[541] ^ message[562] ^ message[563] ^ message[564] ^ message[565] ^ message[566] ^ message[567] ^ message[568] ^ message[569] ^ message[570] ^ message[571] ^ message[572] ^ message[573] ^ message[574] ^ message[575] ^ message[576] ^ message[592] ^ message[593] ^ message[594] ^ message[595] ^ message[596] ^ message[597] ^ message[618] ^ message[619] ^ message[620] ^ message[621] ^ message[622] ^ message[623] ^ message[624] ^ message[625] ^ message[626] ^ message[627] ^ message[628] ^ message[629] ^ message[630] ^ message[631] ^ message[632] ^ message[648] ^ message[649] ^ message[650] ^ message[651] ^ message[652] ^ message[653] ^ message[669] ^ message[670] ^ message[671] ^ message[672] ^ message[673] ^ message[674] ^ message[681] ^ message[697] ^ message[698] ^ message[699] ^ message[700] ^ message[701] ^ message[702] ^ message[703] ^ message[704] ^ message[705] ^ message[706] ^ message[707] ^ message[708] ^ message[709] ^ message[710] ^ message[711] ^ message[712] ^ message[713] ^ message[714] ^ message[715] ^ message[716] ^ message[737] ^ message[738] ^ message[739] ^ message[740] ^ message[741] ^ message[742] ^ message[743] ^ message[744] ^ message[745] ^ message[746] ^ message[747] ^ message[748] ^ message[749] ^ message[750] ^ message[751] ^ message[772] ^ message[773] ^ message[774] ^ message[775] ^ message[776] ^ message[777] ^ message[778] ^ message[779] ^ message[780] ^ message[781] ^ message[782] ^ message[783] ^ message[784] ^ message[785] ^ message[786] ^ message[802] ^ message[803] ^ message[804] ^ message[805] ^ message[806] ^ message[807] ^ message[828] ^ message[829] ^ message[830] ^ message[831] ^ message[832] ^ message[833] ^ message[834] ^ message[835] ^ message[836] ^ message[837] ^ message[838] ^ message[839] ^ message[840] ^ message[841] ^ message[842] ^ message[858] ^ message[859] ^ message[860] ^ message[861] ^ message[862] ^ message[863] ^ message[879] ^ message[880] ^ message[881] ^ message[882] ^ message[883] ^ message[884] ^ message[891] ^ message[912] ^ message[913] ^ message[914] ^ message[915] ^ message[916] ^ message[917] ^ message[918] ^ message[919] ^ message[920] ^ message[921] ^ message[922] ^ message[923] ^ message[924] ^ message[925] ^ message[926] ^ message[942] ^ message[943] ^ message[944] ^ message[945] ^ message[946] ^ message[947] ^ message[963] ^ message[964] ^ message[965] ^ message[966] ^ message[967] ^ message[968] ^ message[975] ^ message[991] ^ message[992] ^ message[993] ^ message[994] ^ message[995] ^ message[996] ^ message[1003] ^ message[1010] ^ message[1012] ^ message[1014] ^ message[1015] ^ message[1016] ^ message[1017] ^ message[1018] ^ message[1019] ^ message[1021] ^ message[1022] ^ message[1023];
    assign parity[6] = message[10] ^ message[11] ^ message[12] ^ message[13] ^ message[14] ^ message[15] ^ message[16] ^ message[17] ^ message[18] ^ message[19] ^ message[30] ^ message[31] ^ message[32] ^ message[33] ^ message[34] ^ message[45] ^ message[46] ^ message[47] ^ message[48] ^ message[49] ^ message[55] ^ message[66] ^ message[67] ^ message[68] ^ message[69] ^ message[70] ^ message[76] ^ message[82] ^ message[94] ^ message[95] ^ message[96] ^ message[97] ^ message[98] ^ message[104] ^ message[110] ^ message[117] ^ message[130] ^ message[131] ^ message[132] ^ message[133] ^ message[134] ^ message[140] ^ message[146] ^ message[153] ^ message[161] ^ message[175] ^ message[176] ^ message[177] ^ message[178] ^ message[179] ^ message[185] ^ message[191] ^ message[198] ^ message[206] ^ message[215] ^ message[221] ^ message[222] ^ message[223] ^ message[224] ^ message[225] ^ message[231] ^ message[232] ^ message[233] ^ message[234] ^ message[235] ^ message[236] ^ message[237] ^ message[238] ^ message[239] ^ message[240] ^ message[246] ^ message[247] ^ message[248] ^ message[249] ^ message[250] ^ message[251] ^ message[252] ^ message[253] ^ message[254] ^ message[255] ^ message[266] ^ message[267] ^ message[268] ^ message[269] ^ message[270] ^ message[271] ^ message[272] ^ message[273] ^ message[274] ^ message[275] ^ message[281] ^ message[282] ^ message[283] ^ message[284] ^ message[285] ^ message[286] ^ message[287] ^ message[288] ^ message[289] ^ message[290] ^ message[301] ^ message[302] ^ message[303] ^ message[304] ^ message[305] ^ message[306] ^ message[307] ^ message[308] ^ message[309] ^ message[310] ^ message[321] ^ message[322] ^ message[323] ^ message[324] ^ message[325] ^ message[326] ^ message[327] ^ message[328] ^ message[329] ^ message[330] ^ message[341] ^ message[342] ^ message[343] ^ message[344] ^ message[345] ^ message[351] ^ message[352] ^ message[353] ^ message[354] ^ message[355] ^ message[356] ^ message[357] ^ message[358] ^ message[359] ^ message[360] ^ message[371] ^ message[372] ^ message[373] ^ message[374] ^ message[375] ^ message[376] ^ message[377] ^ message[378] ^ message[379] ^ message[380] ^ message[391] ^ message[392] ^ message[393] ^ message[394] ^ message[395] ^ message[396] ^ message[397] ^ message[398] ^ message[399] ^ message[400] ^ message[411] ^ message[412] ^ message[413] ^ message[414] ^ message[415] ^ message[426] ^ message[427] ^ message[428] ^ message[429] ^ message[430] ^ message[431] ^ message[432] ^ message[433] ^ message[434] ^ message[435] ^ message[446] ^ message[447] ^ message[448] ^ message[449] ^ message[450] ^ message[461] ^ message[462] ^ message[463] ^ message[464] ^ message[465] ^ message[471] ^ message[477] ^ message[478] ^ message[479] ^ message[480] ^ message[481] ^ message[482] ^ message[483] ^ message[484] ^ message[485] ^ message[486] ^ message[497] ^ message[498] ^ message[499] ^ message[500] ^ message[501] ^ message[502] ^ message[503] ^ message[504] ^ message[505] ^ message[506] ^ message[517] ^ message[518] ^ message[519] ^ message[520] ^ message[521] ^ message[522] ^ message[523] ^ message[524] ^ message[525] ^ message[526] ^ message[537] ^ message[538] ^ message[539] ^ message[540] ^ message[541] ^ message[552] ^ message[553] ^ message[554] ^ message[555] ^ message[556] ^ message[557] ^ message[558] ^ message[559] ^ message[560] ^ message[561] ^ message[572] ^ message[573] ^ message[574] ^ message[575] ^ message[576] ^ message[587] ^ message[588] ^ message[589] ^ message[590] ^ message[591] ^ message[597] ^ message[608] ^ message[609] ^ message[610] ^ message[611] ^ message[612] ^ message[613] ^ message[614] ^ message[615] ^ message[616] ^ message[617] ^ message[628] ^ message[629] ^ message[630] ^ message[631] ^ message[632] ^ message[643] ^ message[644] ^ message[645] ^ message[646] ^ message[647] ^ message[653] ^ message[664] ^ message[665] ^ message[666] ^ message[667] ^ message[668] ^ message[674] ^ message[680] ^ message[687] ^ message[688] ^ message[689] ^ message[690] ^ message[691] ^ message[692] ^ message[693] ^ message[694] ^ message[695] ^ message[696] ^ message[707] ^ message[708] ^ message[709] ^ message[710] ^ message[711] ^ message[712] ^ message[713] ^ message[714] ^ message[715] ^ message[716] ^ message[727] ^ message[728] ^ message[729] ^ message[730] ^ message[731] ^ message[732] ^ message[733] ^ message[734] ^ message[735] ^ message[736] ^ message[747] ^ message[748] ^ message[749] ^ message[750] ^ message[751] ^ message[762] ^ message[763] ^ message[764] ^ message[765] ^ message[766] ^ message[767] ^ message[768] ^ message[769] ^ message[770] ^ message[771] ^ message[782] ^ message[783] ^ message[784] ^ message[785] ^ message[786] ^ message[797] ^ message[798] ^ message[799] ^ message[800] ^ message[801] ^ message[807] ^ message[818] ^ message[819] ^ message[820] ^ message[821] ^ message[822] ^ message[823] ^ message[824] ^ message[825] ^ message[826] ^ message[827] ^ message[838] ^ message[839] ^ message[840] ^ message[841] ^ message[842] ^ message[853] ^ message[854] ^ message[855] ^ message[856] ^ message[857] ^ message[863] ^ message[874] ^ message[875] ^ message[876] ^ message[877] ^ message[878] ^ message[884] ^ message[890] ^ message[902] ^ message[903] ^ message[904] ^ message[905] ^ message[906] ^ message[907] ^ message[908] ^ message[909] ^ message[910] ^ message[911] ^ message[922] ^ message[923] ^ message[924] ^ message[925] ^ message[926] ^ message[937] ^ message[938] ^ message[939] ^ message[940] ^ message[941] ^ message[947] ^ message[958] ^ message[959] ^ message[960] ^ message[961] ^ message[962] ^ message[968] ^ message[974] ^ message[986] ^ message[987] ^ message[988] ^ message[989] ^ message[990] ^ message[996] ^ message[1002] ^ message[1009] ^ message[1012] ^ message[1013] ^ message[1015] ^ message[1016] ^ message[1017] ^ message[1018] ^ message[1019] ^ message[1020] ^ message[1022] ^ message[1023];
    assign parity[7] = message[4] ^ message[5] ^ message[6] ^ message[7] ^ message[8] ^ message[9] ^ message[16] ^ message[17] ^ message[18] ^ message[19] ^ message[26] ^ message[27] ^ message[28] ^ message[29] ^ message[34] ^ message[41] ^ message[42] ^ message[43] ^ message[44] ^ message[49] ^ message[54] ^ message[62] ^ message[63] ^ message[64] ^ message[65] ^ message[70] ^ message[75] ^ message[81] ^ message[90] ^ message[91] ^ message[92] ^ message[93] ^ message[98] ^ message[103] ^ message[109] ^ message[116] ^ message[126] ^ message[127] ^ message[128] ^ message[129] ^ message[134] ^ message[139] ^ message[145] ^ message[152] ^ message[160] ^ message[171] ^ message[172] ^ message[173] ^ message[174] ^ message[179] ^ message[184] ^ message[190] ^ message[197] ^ message[205] ^ message[214] ^ message[220] ^ message[222] ^ message[223] ^ message[224] ^ message[225] ^ message[227] ^ message[228] ^ message[229] ^ message[230] ^ message[235] ^ message[236] ^ message[237] ^ message[238] ^ message[239] ^ message[240] ^ message[242] ^ message[243] ^ message[244] ^ message[245] ^ message[250] ^ message[251] ^ message[252] ^ message[253] ^ message[254] ^ message[255] ^ message[260] ^ message[261] ^ message[262] ^ message[263] ^ message[264] ^ message[265] ^ message[272] ^ message[273] ^ message[274] ^ message[275] ^ message[277] ^ message[278] ^ message[279] ^ message[280] ^ message[285] ^ message[286] ^ message[287] ^ message[288] ^ message[289] ^ message[290] ^ message[295] ^ message[296] ^ message[297] ^ message[298] ^ message[299] ^ message[300] ^ message[307] ^ message[308] ^ message[309] ^ message[310] ^ message[315] ^ message[316] ^ message[317] ^ message[318] ^ message[319] ^ message[320] ^ message[327] ^ message[328] ^ message[329] ^ message[330] ^ message[337] ^ message[338] ^ message[339] ^ message[340] ^ message[345] ^ message[347] ^ message[348] ^ message[349] ^ message[350] ^ message[355] ^ message[356] ^ message[357] ^ message[358] ^ message[359] ^ message[360] ^ message[365] ^ message[366] ^ message[367] ^ message[368] ^ message[369] ^ message[370] ^ message[377] ^ message[378] ^ message[379] ^ message[380] ^ message[385] ^ message[386] ^ message[387] ^ message[388] ^ message[389] ^ message[390] ^ message[397] ^ message[398] ^ message[399] ^ message[400] ^ message[407] ^ message[408] ^ message[409] ^ message[410] ^ message[415] ^ message[420] ^ message[421] ^ message[422] ^ message[423] ^ message[424] ^ message[425] ^ message[432] ^ message[433] ^ message[434] ^ message[435] ^ message[442] ^ message[443] ^ message[444] ^ message[445] ^ message[450] ^ message[457] ^ message[458] ^ message[459] ^ message[460] ^ message[465] ^ message[470] ^ message[473] ^ message[474] ^ message[475] ^ message[476] ^ message[481] ^ message[482] ^ message[483] ^ message[484] ^ message[485] ^ message[486] ^ message[491] ^ message[492] ^ message[493] ^ message[494] ^ message[495] ^ message[496] ^ message[503] ^ message[504] ^ message[505] ^ message[506] ^ message[511] ^ message[512] ^ message[513] ^ message[514] ^ message[515] ^ message[516] ^ message[523] ^ message[524] ^ message[525] ^ message[526] ^ message[533] ^ message[534] ^ message[535] ^ message[536] ^ message[541] ^ message[546] ^ message[547] ^ message[548] ^ message[549] ^ message[550] ^ message[551] ^ message[558] ^ message[559] ^ message[560] ^ message[561] ^ message[568] ^ message[569] ^ message[570] ^ message[571] ^ message[576] ^ message[583] ^ message[584] ^ message[585] ^ message[586] ^ message[591] ^ message[596] ^ message[602] ^ message[603] ^ message[604] ^ message[605] ^ message[606] ^ message[607] ^ message[614] ^ message[615] ^ message[616] ^ message[617] ^ message[624] ^ message[625] ^ message[626] ^ message[627] ^ message[632] ^ message[639] ^ message[640] ^ message[641] ^ message[642] ^ message[647] ^ message[652] ^ message[660] ^ message[661] ^ message[662] ^ message[663] ^ message[668] ^ message[673] ^ message[679] ^ message[683] ^ message[684] ^ message[685] ^ message[686] ^ message[691] ^ message[692] ^ message[693] ^ message[694] ^ message[695] ^ message[696] ^ message[701] ^ message[702] ^ message[703] ^ message[704] ^ message[705] ^ message[706] ^ message[713] ^ message[714] ^ message[715] ^ message[716] ^ message[721] ^ message[722] ^ message[723] ^ message[724] ^ message[725] ^ message[726] ^ message[733] ^ message[734] ^ message[735] ^ message[736] ^ message[743] ^ message[744] ^ message[745] ^ message[746] ^ message[751] ^ message[756] ^ message[757] ^ message[758] ^ message[759] ^ message[760] ^ message[761] ^ message[768] ^ message[769] ^ message[770] ^ message[771] ^ message[778] ^ message[779] ^ message[780] ^ message[781] ^ message[786] ^ message[793] ^ message[794] ^ message[795] ^ message[796] ^ message[801] ^ message[806] ^ message[812] ^ message[813] ^ message[814] ^ message[815] ^ message[816] ^ message[817] ^ message[824] ^ message[825] ^ message[826] ^ message[827] ^ message[834] ^ message[835] ^ message[836] ^ message[837] ^ message[842] ^ message[849] ^ message[850] ^ message[851] ^ message[852] ^ message[857] ^ message[862] ^ message[870] ^ message[871] ^ message[872] ^ message[873] ^ message[878] ^ message[883] ^ message[889] ^ message[896] ^ message[897] ^ message[898] ^ message[899] ^ message[900] ^ message[901] ^ message[908] ^ message[909] ^ message[910] ^ message[911] ^ message[918] ^ message[919] ^ message[920] ^ message[921] ^ message[926] ^ message[933] ^ message[934] ^ message[935] ^ message[936] ^ message[941] ^ message[946] ^ message[954] ^ message[955] ^ message[956] ^ message[957] ^ message[962] ^ message[967] ^ message[973] ^ message[982] ^ message[983] ^ message[984] ^ message[985] ^ message[990] ^ message[995] ^ message[1001] ^ message[1008] ^ message[1012] ^ message[1013] ^ message[1014] ^ message[1016] ^ message[1017] ^ message[1018] ^ message[1019] ^ message[1020] ^ message[1021] ^ message[1023];
    assign parity[8] = message[1] ^ message[2] ^ message[3] ^ message[7] ^ message[8] ^ message[9] ^ message[13] ^ message[14] ^ message[15] ^ message[19] ^ message[23] ^ message[24] ^ message[25] ^ message[29] ^ message[33] ^ message[38] ^ message[39] ^ message[40] ^ message[44] ^ message[48] ^ message[53] ^ message[59] ^ message[60] ^ message[61] ^ message[65] ^ message[69] ^ message[74] ^ message[80] ^ message[87] ^ message[88] ^ message[89] ^ message[93] ^ message[97] ^ message[102] ^ message[108] ^ message[115] ^ message[123] ^ message[124] ^ message[125] ^ message[129] ^ message[133] ^ message[138] ^ message[144] ^ message[151] ^ message[159] ^ message[168] ^ message[169] ^ message[170] ^ message[174] ^ message[178] ^ message[183] ^ message[189] ^ message[196] ^ message[204] ^ message[213] ^ message[220] ^ message[221] ^ message[223] ^ message[224] ^ message[225] ^ message[226] ^ message[228] ^ message[229] ^ message[230] ^ message[232] ^ message[233] ^ message[234] ^ message[238] ^ message[239] ^ message[240] ^ message[241] ^ message[243] ^ message[244] ^ message[245] ^ message[247] ^ message[248] ^ message[249] ^ message[253] ^ message[254] ^ message[255] ^ message[257] ^ message[258] ^ message[259] ^ message[263] ^ message[264] ^ message[265] ^ message[269] ^ message[270] ^ message[271] ^ message[275] ^ message[276] ^ message[278] ^ message[279] ^ message[280] ^ message[282] ^ message[283] ^ message[284] ^ message[288] ^ message[289] ^ message[290] ^ message[292] ^ message[293] ^ message[294] ^ message[298] ^ message[299] ^ message[300] ^ message[304] ^ message[305] ^ message[306] ^ message[310] ^ message[312] ^ message[313] ^ message[314] ^ message[318] ^ message[319] ^ message[320] ^ message[324] ^ message[325] ^ message[326] ^ message[330] ^ message[334] ^ message[335] ^ message[336] ^ message[340] ^ message[344] ^ message[346] ^ message[348] ^ message[349] ^ message[350] ^ message[352] ^ message[353] ^ message[354] ^ message[358] ^ message[359] ^ message[360] ^ message[362] ^ message[363] ^ message[364] ^ message[368] ^ message[369] ^ message[370] ^ message[374] ^ message[375] ^ message[376] ^ message[380] ^ message[382] ^ message[383] ^ message[384] ^ message[388] ^ message[389] ^ message[390] ^ message[394] ^ message[395] ^ message[396] ^ message[400] ^ message[404] ^ message[405] ^ message[406] ^ message[410] ^ message[414] ^ message[417] ^ message[418] ^ message[419] ^ message[423] ^ message[424] ^ message[425] ^ message[429] ^ message[430] ^ message[431] ^ message[435] ^ message[439] ^ message[440] ^ message[441] ^ message[445] ^ message[449] ^ message[454] ^ message[455] ^ message[456] ^ message[460] ^ message[464] ^ message[469] ^ message[472] ^ message[474] ^ message[475] ^ message[476] ^ message[478] ^ message[479] ^ message[480] ^ message[484] ^ message[485] ^ message[486] ^ message[488] ^ message[489] ^ message[490] ^ message[494] ^ message[495] ^ message[496] ^ message[500] ^ message[501] ^ message[502] ^ message[506] ^ message[508] ^ message[509] ^ message[510] ^ message[514] ^ message[515] ^ message[516] ^ message[520] ^ message[521] ^ message[522] ^ message[526] ^ message[530] ^ message[531] ^ message[532] ^ message[536] ^ message[540] ^ message[543] ^ message[544] ^ message[545] ^ message[549] ^ message[550] ^ message[551] ^ message[555] ^ message[556] ^ message[557] ^ message[561] ^ message[565] ^ message[566] ^ message[567] ^ message[571] ^ message[575] ^ message[580] ^ message[581] ^ message[582] ^ message[586] ^ message[590] ^ message[595] ^ message[599] ^ message[600] ^ message[601] ^ message[605] ^ message[606] ^ message[607] ^ message[611] ^ message[612] ^ message[613] ^ message[617] ^ message[621] ^ message[622] ^ message[623] ^ message[627] ^ message[631] ^ message[636] ^ message[637] ^ message[638] ^ message[642] ^ message[646] ^ message[651] ^ message[657] ^ message[658] ^ message[659] ^ message[663] ^ message[667] ^ message[672] ^ message[678] ^ message[682] ^ message[684] ^ message[685] ^ message[686] ^ message[688] ^ message[689] ^ message[690] ^ message[694] ^ message[695] ^ message[696] ^ message[698] ^ message[699] ^ message[700] ^ message[704] ^ message[705] ^ message[706] ^ message[710] ^ message[711] ^ message[712] ^ message[716] ^ message[718] ^ message[719] ^ message[720] ^ message[724] ^ message[725] ^ message[726] ^ message[730] ^ message[731] ^ message[732] ^ message[736] ^ message[740] ^ message[741] ^ message[742] ^ message[746] ^ message[750] ^ message[753] ^ message[754] ^ message[755] ^ message[759] ^ message[760] ^ message[761] ^ message[765] ^ message[766] ^ message[767] ^ message[771] ^ message[775] ^ message[776] ^ message[777] ^ message[781] ^ message[785] ^ message[790] ^ message[791] ^ message[792] ^ message[796] ^ message[800] ^ message[805] ^ message[809] ^ message[810] ^ message[811] ^ message[815] ^ message[816] ^ message[817] ^ message[821] ^ message[822] ^ message[823] ^ message[827] ^ message[831] ^ message[832] ^ message[833] ^ message[837] ^ message[841] ^ message[846] ^ message[847] ^ message[848] ^ message[852] ^ message[856] ^ message[861] ^ message[867] ^ message[868] ^ message[869] ^ message[873] ^ message[877] ^ message[882] ^ message[888] ^ message[893] ^ message[894] ^ message[895] ^ message[899] ^ message[900] ^ message[901] ^ message[905] ^ message[906] ^ message[907] ^ message[911] ^ message[915] ^ message[916] ^ message[917] ^ message[921] ^ message[925] ^ message[930] ^ message[931] ^ message[932] ^ message[936] ^ message[940] ^ message[945] ^ message[951] ^ message[952] ^ message[953] ^ message[957] ^ message[961] ^ message[966] ^ message[972] ^ message[979] ^ message[980] ^ message[981] ^ message[985] ^ message[989] ^ message[994] ^ message[1000] ^ message[1007] ^ message[1012] ^ message[1013] ^ message[1014] ^ message[1015] ^ message[1017] ^ message[1018] ^ message[1019] ^ message[1020] ^ message[1021] ^ message[1022];
    assign parity[9] = message[0] ^ message[2] ^ message[3] ^ message[5] ^ message[6] ^ message[9] ^ message[11] ^ message[12] ^ message[15] ^ message[18] ^ message[21] ^ message[22] ^ message[25] ^ message[28] ^ message[32] ^ message[36] ^ message[37] ^ message[40] ^ message[43] ^ message[47] ^ message[52] ^ message[57] ^ message[58] ^ message[61] ^ message[64] ^ message[68] ^ message[73] ^ message[79] ^ message[85] ^ message[86] ^ message[89] ^ message[92] ^ message[96] ^ message[101] ^ message[107] ^ message[114] ^ message[121] ^ message[122] ^ message[125] ^ message[128] ^ message[132] ^ message[137] ^ message[143] ^ message[150] ^ message[158] ^ message[166] ^ message[167] ^ message[170] ^ message[173] ^ message[177] ^ message[182] ^ message[188] ^ message[195] ^ message[203] ^ message[212] ^ message[220] ^ message[221] ^ message[222] ^ message[224] ^ message[225] ^ message[226] ^ message[227] ^ message[229] ^ message[230] ^ message[231] ^ message[233] ^ message[234] ^ message[236] ^ message[237] ^ message[240] ^ message[241] ^ message[242] ^ message[244] ^ message[245] ^ message[246] ^ message[248] ^ message[249] ^ message[251] ^ message[252] ^ message[255] ^ message[256] ^ message[258] ^ message[259] ^ message[261] ^ message[262] ^ message[265] ^ message[267] ^ message[268] ^ message[271] ^ message[274] ^ message[276] ^ message[277] ^ message[279] ^ message[280] ^ message[281] ^ message[283] ^ message[284] ^ message[286] ^ message[287] ^ message[290] ^ message[291] ^ message[293] ^ message[294] ^ message[296] ^ message[297] ^ message[300] ^ message[302] ^ message[303] ^ message[306] ^ message[309] ^ message[311] ^ message[313] ^ message[314] ^ message[316] ^ message[317] ^ message[320] ^ message[322] ^ message[323] ^ message[326] ^ message[329] ^ message[332] ^ message[333] ^ message[336] ^ message[339] ^ message[343] ^ message[346] ^ message[347] ^ message[349] ^ message[350] ^ message[351] ^ message[353] ^ message[354] ^ message[356] ^ message[357] ^ message[360] ^ message[361] ^ message[363] ^ message[364] ^ message[366] ^ message[367] ^ message[370] ^ message[372] ^ message[373] ^ message[376] ^ message[379] ^ message[381] ^ message[383] ^ message[384] ^ message[386] ^ message[387] ^ message[390] ^ message[392] ^ message[393] ^ message[396] ^ message[399] ^ message[402] ^ message[403] ^ message[406] ^ message[409] ^ message[413] ^ message[416] ^ message[418] ^ message[419] ^ message[421] ^ message[422] ^ message[425] ^ message[427] ^ message[428] ^ message[431] ^ message[434] ^ message[437] ^ message[438] ^ message[441] ^ message[444] ^ message[448] ^ message[452] ^ message[453] ^ message[456] ^ message[459] ^ message[463] ^ message[468] ^ message[472] ^ message[473] ^ message[475] ^ message[476] ^ message[477] ^ message[479] ^ message[480] ^ message[482] ^ message[483] ^ message[486] ^ message[487] ^ message[489] ^ message[490] ^ message[492] ^ message[493] ^ message[496] ^ message[498] ^ message[499] ^ message[502] ^ message[505] ^ message[507] ^ message[509] ^ message[510] ^ message[512] ^ message[513] ^ message[516] ^ message[518] ^ message[519] ^ message[522] ^ message[525] ^ message[528] ^ message[529] ^ message[532] ^ message[535] ^ message[539] ^ message[542] ^ message[544] ^ message[545] ^ message[547] ^ message[548] ^ message[551] ^ message[553] ^ message[554] ^ message[557] ^ message[560] ^ message[563] ^ message[564] ^ message[567] ^ message[570] ^ message[574] ^ message[578] ^ message[579] ^ message[582] ^ message[585] ^ message[589] ^ message[594] ^ message[598] ^ message[600] ^ message[601] ^ message[603] ^ message[604] ^ message[607] ^ message[609] ^ message[610] ^ message[613] ^ message[616] ^ message[619] ^ message[620] ^ message[623] ^ message[626] ^ message[630] ^ message[634] ^ message[635] ^ message[638] ^ message[641] ^ message[645] ^ message[650] ^ message[655] ^ message[656] ^ message[659] ^ message[662] ^ message[666] ^ message[671] ^ message[677] ^ message[682] ^ message[683] ^ message[685] ^ message[686] ^ message[687] ^ message[689] ^ message[690] ^ message[692] ^ message[693] ^ message[696] ^ message[697] ^ message[699] ^ message[700] ^ message[702] ^ message[703] ^ message[706] ^ message[708] ^ message[709] ^ message[712] ^ message[715] ^ message[717] ^ message[719] ^ message[720] ^ message[722] ^ message[723] ^ message[726] ^ message[728] ^ message[729] ^ message[732] ^ message[735] ^ message[738] ^ message[739] ^ message[742] ^ message[745] ^ message[749] ^ message[752] ^ message[754] ^ message[755] ^ message[757] ^ message[758] ^ message[761] ^ message[763] ^ message[764] ^ message[767] ^ message[770] ^ message[773] ^ message[774] ^ message[777] ^ message[780] ^ message[784] ^ message[788] ^ message[789] ^ message[792] ^ message[795] ^ message[799] ^ message[804] ^ message[808] ^ message[810] ^ message[811] ^ message[813] ^ message[814] ^ message[817] ^ message[819] ^ message[820] ^ message[823] ^ message[826] ^ message[829] ^ message[830] ^ message[833] ^ message[836] ^ message[840] ^ message[844] ^ message[845] ^ message[848] ^ message[851] ^ message[855] ^ message[860] ^ message[865] ^ message[866] ^ message[869] ^ message[872] ^ message[876] ^ message[881] ^ message[887] ^ message[892] ^ message[894] ^ message[895] ^ message[897] ^ message[898] ^ message[901] ^ message[903] ^ message[904] ^ message[907] ^ message[910] ^ message[913] ^ message[914] ^ message[917] ^ message[920] ^ message[924] ^ message[928] ^ message[929] ^ message[932] ^ message[935] ^ message[939] ^ message[944] ^ message[949] ^ message[950] ^ message[953] ^ message[956] ^ message[960] ^ message[965] ^ message[971] ^ message[977] ^ message[978] ^ message[981] ^ message[984] ^ message[988] ^ message[993] ^ message[999] ^ message[1006] ^ message[1012] ^ message[1013] ^ message[1014] ^ message[1015] ^ message[1016] ^ message[1018] ^ message[1019] ^ message[1020] ^ message[1021] ^ message[1022] ^ message[1023];
    assign parity[10] = message[0] ^ message[1] ^ message[3] ^ message[4] ^ message[6] ^ message[8] ^ message[10] ^ message[12] ^ message[14] ^ message[17] ^ message[20] ^ message[22] ^ message[24] ^ message[27] ^ message[31] ^ message[35] ^ message[37] ^ message[39] ^ message[42] ^ message[46] ^ message[51] ^ message[56] ^ message[58] ^ message[60] ^ message[63] ^ message[67] ^ message[72] ^ message[78] ^ message[84] ^ message[86] ^ message[88] ^ message[91] ^ message[95] ^ message[100] ^ message[106] ^ message[113] ^ message[120] ^ message[122] ^ message[124] ^ message[127] ^ message[131] ^ message[136] ^ message[142] ^ message[149] ^ message[157] ^ message[165] ^ message[167] ^ message[169] ^ message[172] ^ message[176] ^ message[181] ^ message[187] ^ message[194] ^ message[202] ^ message[211] ^ message[220] ^ message[221] ^ message[222] ^ message[223] ^ message[225] ^ message[226] ^ message[227] ^ message[228] ^ message[230] ^ message[231] ^ message[232] ^ message[234] ^ message[235] ^ message[237] ^ message[239] ^ message[241] ^ message[242] ^ message[243] ^ message[245] ^ message[246] ^ message[247] ^ message[249] ^ message[250] ^ message[252] ^ message[254] ^ message[256] ^ message[257] ^ message[259] ^ message[260] ^ message[262] ^ message[264] ^ message[266] ^ message[268] ^ message[270] ^ message[273] ^ message[276] ^ message[277] ^ message[278] ^ message[280] ^ message[281] ^ message[282] ^ message[284] ^ message[285] ^ message[287] ^ message[289] ^ message[291] ^ message[292] ^ message[294] ^ message[295] ^ message[297] ^ message[299] ^ message[301] ^ message[303] ^ message[305] ^ message[308] ^ message[311] ^ message[312] ^ message[314] ^ message[315] ^ message[317] ^ message[319] ^ message[321] ^ message[323] ^ message[325] ^ message[328] ^ message[331] ^ message[333] ^ message[335] ^ message[338] ^ message[342] ^ message[346] ^ message[347] ^ message[348] ^ message[350] ^ message[351] ^ message[352] ^ message[354] ^ message[355] ^ message[357] ^ message[359] ^ message[361] ^ message[362] ^ message[364] ^ message[365] ^ message[367] ^ message[369] ^ message[371] ^ message[373] ^ message[375] ^ message[378] ^ message[381] ^ message[382] ^ message[384] ^ message[385] ^ message[387] ^ message[389] ^ message[391] ^ message[393] ^ message[395] ^ message[398] ^ message[401] ^ message[403] ^ message[405] ^ message[408] ^ message[412] ^ message[416] ^ message[417] ^ message[419] ^ message[420] ^ message[422] ^ message[424] ^ message[426] ^ message[428] ^ message[430] ^ message[433] ^ message[436] ^ message[438] ^ message[440] ^ message[443] ^ message[447] ^ message[451] ^ message[453] ^ message[455] ^ message[458] ^ message[462] ^ message[467] ^ message[472] ^ message[473] ^ message[474] ^ message[476] ^ message[477] ^ message[478] ^ message[480] ^ message[481] ^ message[483] ^ message[485] ^ message[487] ^ message[488] ^ message[490] ^ message[491] ^ message[493] ^ message[495] ^ message[497] ^ message[499] ^ message[501] ^ message[504] ^ message[507] ^ message[508] ^ message[510] ^ message[511] ^ message[513] ^ message[515] ^ message[517] ^ message[519] ^ message[521] ^ message[524] ^ message[527] ^ message[529] ^ message[531] ^ message[534] ^ message[538] ^ message[542] ^ message[543] ^ message[545] ^ message[546] ^ message[548] ^ message[550] ^ message[552] ^ message[554] ^ message[556] ^ message[559] ^ message[562] ^ message[564] ^ message[566] ^ message[569] ^ message[573] ^ message[577] ^ message[579] ^ message[581] ^ message[584] ^ message[588] ^ message[593] ^ message[598] ^ message[599] ^ message[601] ^ message[602] ^ message[604] ^ message[606] ^ message[608] ^ message[610] ^ message[612] ^ message[615] ^ message[618] ^ message[620] ^ message[622] ^ message[625] ^ message[629] ^ message[633] ^ message[635] ^ message[637] ^ message[640] ^ message[644] ^ message[649] ^ message[654] ^ message[656] ^ message[658] ^ message[661] ^ message[665] ^ message[670] ^ message[676] ^ message[682] ^ message[683] ^ message[684] ^ message[686] ^ message[687] ^ message[688] ^ message[690] ^ message[691] ^ message[693] ^ message[695] ^ message[697] ^ message[698] ^ message[700] ^ message[701] ^ message[703] ^ message[705] ^ message[707] ^ message[709] ^ message[711] ^ message[714] ^ message[717] ^ message[718] ^ message[720] ^ message[721] ^ message[723] ^ message[725] ^ message[727] ^ message[729] ^ message[731] ^ message[734] ^ message[737] ^ message[739] ^ message[741] ^ message[744] ^ message[748] ^ message[752] ^ message[753] ^ message[755] ^ message[756] ^ message[758] ^ message[760] ^ message[762] ^ message[764] ^ message[766] ^ message[769] ^ message[772] ^ message[774] ^ message[776] ^ message[779] ^ message[783] ^ message[787] ^ message[789] ^ message[791] ^ message[794] ^ message[798] ^ message[803] ^ message[808] ^ message[809] ^ message[811] ^ message[812] ^ message[814] ^ message[816] ^ message[818] ^ message[820] ^ message[822] ^ message[825] ^ message[828] ^ message[830] ^ message[832] ^ message[835] ^ message[839] ^ message[843] ^ message[845] ^ message[847] ^ message[850] ^ message[854] ^ message[859] ^ message[864] ^ message[866] ^ message[868] ^ message[871] ^ message[875] ^ message[880] ^ message[886] ^ message[892] ^ message[893] ^ message[895] ^ message[896] ^ message[898] ^ message[900] ^ message[902] ^ message[904] ^ message[906] ^ message[909] ^ message[912] ^ message[914] ^ message[916] ^ message[919] ^ message[923] ^ message[927] ^ message[929] ^ message[931] ^ message[934] ^ message[938] ^ message[943] ^ message[948] ^ message[950] ^ message[952] ^ message[955] ^ message[959] ^ message[964] ^ message[970] ^ message[976] ^ message[978] ^ message[980] ^ message[983] ^ message[987] ^ message[992] ^ message[998] ^ message[1005] ^ message[1012] ^ message[1013] ^ message[1014] ^ message[1015] ^ message[1016] ^ message[1017] ^ message[1019] ^ message[1020] ^ message[1021] ^ message[1022] ^ message[1023];
    assign parity[11] = message[0] ^ message[1] ^ message[2] ^ message[4] ^ message[5] ^ message[7] ^ message[10] ^ message[11] ^ message[13] ^ message[16] ^ message[20] ^ message[21] ^ message[23] ^ message[26] ^ message[30] ^ message[35] ^ message[36] ^ message[38] ^ message[41] ^ message[45] ^ message[50] ^ message[56] ^ message[57] ^ message[59] ^ message[62] ^ message[66] ^ message[71] ^ message[77] ^ message[84] ^ message[85] ^ message[87] ^ message[90] ^ message[94] ^ message[99] ^ message[105] ^ message[112] ^ message[120] ^ message[121] ^ message[123] ^ message[126] ^ message[130] ^ message[135] ^ message[141] ^ message[148] ^ message[156] ^ message[165] ^ message[166] ^ message[168] ^ message[171] ^ message[175] ^ message[180] ^ message[186] ^ message[193] ^ message[201] ^ message[210] ^ message[220] ^ message[221] ^ message[222] ^ message[223] ^ message[224] ^ message[226] ^ message[227] ^ message[228] ^ message[229] ^ message[231] ^ message[232] ^ message[233] ^ message[235] ^ message[236] ^ message[238] ^ message[241] ^ message[242] ^ message[243] ^ message[244] ^ message[246] ^ message[247] ^ message[248] ^ message[250] ^ message[251] ^ message[253] ^ message[256] ^ message[257] ^ message[258] ^ message[260] ^ message[261] ^ message[263] ^ message[266] ^ message[267] ^ message[269] ^ message[272] ^ message[276] ^ message[277] ^ message[278] ^ message[279] ^ message[281] ^ message[282] ^ message[283] ^ message[285] ^ message[286] ^ message[288] ^ message[291] ^ message[292] ^ message[293] ^ message[295] ^ message[296] ^ message[298] ^ message[301] ^ message[302] ^ message[304] ^ message[307] ^ message[311] ^ message[312] ^ message[313] ^ message[315] ^ message[316] ^ message[318] ^ message[321] ^ message[322] ^ message[324] ^ message[327] ^ message[331] ^ message[332] ^ message[334] ^ message[337] ^ message[341] ^ message[346] ^ message[347] ^ message[348] ^ message[349] ^ message[351] ^ message[352] ^ message[353] ^ message[355] ^ message[356] ^ message[358] ^ message[361] ^ message[362] ^ message[363] ^ message[365] ^ message[366] ^ message[368] ^ message[371] ^ message[372] ^ message[374] ^ message[377] ^ message[381] ^ message[382] ^ message[383] ^ message[385] ^ message[386] ^ message[388] ^ message[391] ^ message[392] ^ message[394] ^ message[397] ^ message[401] ^ message[402] ^ message[404] ^ message[407] ^ message[411] ^ message[416] ^ message[417] ^ message[418] ^ message[420] ^ message[421] ^ message[423] ^ message[426] ^ message[427] ^ message[429] ^ message[432] ^ message[436] ^ message[437] ^ message[439] ^ message[442] ^ message[446] ^ message[451] ^ message[452] ^ message[454] ^ message[457] ^ message[461] ^ message[466] ^ message[472] ^ message[473] ^ message[474] ^ message[475] ^ message[477] ^ message[478] ^ message[479] ^ message[481] ^ message[482] ^ message[484] ^ message[487] ^ message[488] ^ message[489] ^ message[491] ^ message[492] ^ message[494] ^ message[497] ^ message[498] ^ message[500] ^ message[503] ^ message[507] ^ message[508] ^ message[509] ^ message[511] ^ message[512] ^ message[514] ^ message[517] ^ message[518] ^ message[520] ^ message[523] ^ message[527] ^ message[528] ^ message[530] ^ message[533] ^ message[537] ^ message[542] ^ message[543] ^ message[544] ^ message[546] ^ message[547] ^ message[549] ^ message[552] ^ message[553] ^ message[555] ^ message[558] ^ message[562] ^ message[563] ^ message[565] ^ message[568] ^ message[572] ^ message[577] ^ message[578] ^ message[580] ^ message[583] ^ message[587] ^ message[592] ^ message[598] ^ message[599] ^ message[600] ^ message[602] ^ message[603] ^ message[605] ^ message[608] ^ message[609] ^ message[611] ^ message[614] ^ message[618] ^ message[619] ^ message[621] ^ message[624] ^ message[628] ^ message[633] ^ message[634] ^ message[636] ^ message[639] ^ message[643] ^ message[648] ^ message[654] ^ message[655] ^ message[657] ^ message[660] ^ message[664] ^ message[669] ^ message[675] ^ message[682] ^ message[683] ^ message[684] ^ message[685] ^ message[687] ^ message[688] ^ message[689] ^ message[691] ^ message[692] ^ message[694] ^ message[697] ^ message[698] ^ message[699] ^ message[701] ^ message[702] ^ message[704] ^ message[707] ^ message[708] ^ message[710] ^ message[713] ^ message[717] ^ message[718] ^ message[719] ^ message[721] ^ message[722] ^ message[724] ^ message[727] ^ message[728] ^ message[730] ^ message[733] ^ message[737] ^ message[738] ^ message[740] ^ message[743] ^ message[747] ^ message[752] ^ message[753] ^ message[754] ^ message[756] ^ message[757] ^ message[759] ^ message[762] ^ message[763] ^ message[765] ^ message[768] ^ message[772] ^ message[773] ^ message[775] ^ message[778] ^ message[782] ^ message[787] ^ message[788] ^ message[790] ^ message[793] ^ message[797] ^ message[802] ^ message[808] ^ message[809] ^ message[810] ^ message[812] ^ message[813] ^ message[815] ^ message[818] ^ message[819] ^ message[821] ^ message[824] ^ message[828] ^ message[829] ^ message[831] ^ message[834] ^ message[838] ^ message[843] ^ message[844] ^ message[846] ^ message[849] ^ message[853] ^ message[858] ^ message[864] ^ message[865] ^ message[867] ^ message[870] ^ message[874] ^ message[879] ^ message[885] ^ message[892] ^ message[893] ^ message[894] ^ message[896] ^ message[897] ^ message[899] ^ message[902] ^ message[903] ^ message[905] ^ message[908] ^ message[912] ^ message[913] ^ message[915] ^ message[918] ^ message[922] ^ message[927] ^ message[928] ^ message[930] ^ message[933] ^ message[937] ^ message[942] ^ message[948] ^ message[949] ^ message[951] ^ message[954] ^ message[958] ^ message[963] ^ message[969] ^ message[976] ^ message[977] ^ message[979] ^ message[982] ^ message[986] ^ message[991] ^ message[997] ^ message[1004] ^ message[1012] ^ message[1013] ^ message[1014] ^ message[1015] ^ message[1016] ^ message[1017] ^ message[1018] ^ message[1020] ^ message[1021] ^ message[1022] ^ message[1023];
  end else begin : gen_default_parity
    `BR_ASSERT_STATIC(invalid_parity_width_a, 1'b0)
  end

  // ri lint_check_on EXPR_ID_LIMIT

  //------
  // Concatenate message and parity bits to form the codeword.
  //------
  logic [CodewordWidth-1:0] internal_codeword;
  assign internal_codeword = {parity, message};

  //------
  // Optionally register the output signals.
  //------
  br_delay_valid #(
      .Width(CodewordWidth),
      .NumStages(RegisterOutputs == 1 ? 1 : 0)
  ) br_delay_valid_outputs (
      .clk,
      .rst,
      .in_valid(data_valid),
      .in({internal_codeword}),
      .out_valid(codeword_valid),
      .out(codeword),
      .out_valid_stages(),  // unused
      .out_stages()  // unused
  );

  //------------------------------------------
  // Implementation checks
  //------------------------------------------
  `BR_ASSERT_IMPL(latency_a, data_valid |-> ##Latency codeword_valid)

  // verilog_lint: waive-stop line-length
  // verilog_format: on

endmodule : br_ecc_secded_encoder
