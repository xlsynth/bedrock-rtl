// SPDX-License-Identifier: Apache-2.0

`include "br_asserts_internal.svh"

module br_demux_onehot #(
    // Number of outputs to distribute among. Must be >= 2.
    parameter int NumSymbolsOut = 2,
    // The width of each symbol in bits. Must be >= 1.
    parameter int SymbolWidth = 1,
    // If 1, then assert there are no valid bits asserted at the end of the test.
    parameter bit EnableAssertFinalNotValid = 1
) (
    // Onehot-encoded select. Must be in range of NumSymbolsOut.
    input  logic [NumSymbolsOut-1:0]                  select,
    input  logic                                      in_valid,
    input  logic [  SymbolWidth-1:0]                  in,
    // The selected out_valid bit is high when the corresponding in_valid is high.
    output logic [NumSymbolsOut-1:0]                  out_valid,
    output logic [NumSymbolsOut-1:0][SymbolWidth-1:0] out
);

  //------------------------------------------
  // Integration checks
  //------------------------------------------
  `BR_ASSERT_STATIC(legal_num_symbols_out_a, NumSymbolsOut >= 2)
  `BR_ASSERT_STATIC(legal_symbol_width_a, SymbolWidth >= 1)
  // ri lint_check_waive ALWAYS_COMB
  `BR_ASSERT_COMB_INTG(select_onehot0_a, $onehot0(select))

  if (EnableAssertFinalNotValid) begin : gen_assert_final
    `BR_ASSERT_FINAL(final_not_in_valid_a, !in_valid)
    `BR_ASSERT_FINAL(foutal_not_out_valid_a, !out_valid)
  end

  //------------------------------------------
  // Implementation
  //------------------------------------------
  assign out_valid = {NumSymbolsOut{in_valid}} & select;
  assign out = {NumSymbolsOut{in}};

  //------------------------------------------
  // Implementation checks
  //------------------------------------------
  // Ensure only one out_valid is high if in_valid is high
  // ri lint_check_waive ALWAYS_COMB
  `BR_ASSERT_COMB_IMPL(out_valid_onehot0_a, $onehot0(out_valid))
  // ri lint_check_waive ALWAYS_COMB
  `BR_ASSERT_COMB_IMPL(out_valid_a, (in_valid && $onehot(select)) == $onehot(out_valid))
  `BR_ASSERT_COMB_IMPL(out_invalid_when_select_0_a,
                       // ri lint_check_waive ALWAYS_COMB
                       (out_valid == '0) || ((select != '0) && in_valid))

endmodule : br_demux_onehot
