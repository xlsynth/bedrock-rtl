// Copyright 2025 The Bedrock-RTL Authors
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//     http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.

// Bedrock-RTL Delay Line Deskew (Valid-Next to Valid)
//
// Retimes a delay line using skewed valid-next/data (i.e., valid runs one
// cycle ahead of data)to instead use aligned valid/data). Registers the valid while
// letting the data pass through. This is not considered to add datapath latency
// because the incoming valid was already ahead of the data by 1 cycle.
//
// This module has no reset. The valid register will flush from the input.

`include "br_registers.svh"
`include "br_asserts_internal.svh"

module br_delay_deskew #(
    parameter int Width = 1,  // Must be at least 1
    // If 1, then assert there are no valid bits asserted at the end of the test.
    parameter bit EnableAssertFinalNotValid = 1
) (
    // Positive edge-triggered clock.
    input  logic             clk,
    input  logic             in_valid_next,
    input  logic [Width-1:0] in,
    output logic             out_valid,
    output logic [Width-1:0] out
);

  //------------------------------------------
  // Integration checks
  //------------------------------------------
  `BR_ASSERT_STATIC(width_must_be_at_least_one_a, Width >= 1)

  // ri lint_check_waive ALWAYS_COMB
  `BR_COVER_COMB_INTG(in_valid_next_c, in_valid_next)

  if (EnableAssertFinalNotValid) begin : gen_assert_final
    `BR_ASSERT_FINAL(final_not_in_valid_next_a, !in_valid_next)
    `BR_ASSERT_FINAL(final_not_out_valid_a, !out_valid)
  end

  //------------------------------------------
  // Implementation
  //------------------------------------------
  `BR_REGN(out_valid, in_valid_next)
  assign out = in;

  //------------------------------------------
  // Implementation checks
  //------------------------------------------
  `BR_ASSERT_CR_IMPL(valid_delay_a, ##1 out_valid === $past(in_valid_next), clk, 1'b0)
  // ri lint_check_waive ALWAYS_COMB
  `BR_ASSERT_COMB_IMPL(data_delay_a, out === in)

endmodule : br_delay_deskew
