// Copyright 2024-2025 The Bedrock-RTL Authors
//
// Licensed under the Apache License, Version 2.0 (the "License");
// Copyright 2024-2025 The Bedrock-RTL Authors
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//     http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.


// verilog_format: off
// verilog_lint: waive-start line-length

// Bedrock-RTL Single-Error-Correcting, Double-Error-Detecting (SECDED - Hsiao) Decoder
//
// Decodes a codeword using a single-error-correcting, double-error-detecting
// linear block code in systematic form (in layperson's terms: a Hsiao SECDED [1] decoder,
// closely related to Hamming codes).
//
// Systematic form means that the codeword is formed by appending the
// calculated parity bits to the message, i.e., the code has the property
// that the message bits are 1:1 with a slice of bits in the codeword (if they
// have not been corrupted).
//
// In Bedrock ECC libs, our convention is to always append the parity bits on
// the MSbs:
//     codeword == {parity, message}
//
// The data is still marked valid even if an error is detected.
//
// This module has parameterizable latency. By default, it is purely combinational,
// but it can have up to 3 cycles of delay (RegisterInputs, RegisterSyndrome, and
// RegisterOutputs). The initiation interval is always 1 cycle.
//
// Any data width >= 4 is supported, up to a maximum of 1024. It is considered
// internally zero-padded up to the largest message width supported by the number of parity bits
// as part of decoding. The following table outlines the number of parity bits required for
// different message widths.
//
// | Message Width (k) | Parity Width (r) | Codeword Width (n)|
// |-------------------|------------------|-------------------|
// | 4                 | 4                | 8                 |
// | 11                | 5                | 16                |
// | 26                | 6                | 32                |
// | 57                | 7                | 64                |
// | 120               | 8                | 128               |
// | 247               | 9                | 256               |
// | 502               | 10               | 512               |
// | 1013              | 11               | 1024              |
// | 2036              | 12               | 2048              |
//
// The number of parity bits must be one of the values in the table above
// or the module will not elaborate.
//
// References:
// [1] https://ieeexplore.ieee.org/abstract/document/5391627

`include "br_asserts.svh"
`include "br_asserts_internal.svh"
`include "br_assign.svh"
`include "br_unused.svh"

// TODO(mgottscho): Pipeline the syndrome decoding and then correction with a parameter.
module br_ecc_secded_decoder #(
    parameter int DataWidth = 4,  // Must be at least 4
    parameter int ParityWidth = 4,  // Must be at least 4 and at most 12
    // If 1, then insert a pipeline register at the input.
    parameter bit RegisterInputs = 0,
    // If 1, then insert a pipeline register between syndrome computation and
    // syndrome decoding (error correction).
    parameter bit RegisterSyndrome = 0,
    // If 1, then insert a pipeline register at the output.
    parameter bit RegisterOutputs = 0,
    // If 1, then assert there are no valid bits asserted at the end of the test.
    parameter bit EnableAssertFinalNotValid = 1,
    localparam int InputWidth = DataWidth + ParityWidth,
    localparam int MessageWidth = br_ecc::get_max_message_width(ParityWidth),
    localparam int CodewordWidth = MessageWidth + ParityWidth,
    // ri lint_check_waive PARAM_NOT_USED
    localparam int Latency = RegisterInputs + RegisterSyndrome + RegisterOutputs
) (
    // Positive edge-triggered clock.
    input  logic                     clk,
    // Synchronous active-high reset.
    input  logic                     rst,

    // Decoder input (received data and parity, possibly with errors).
    // Provide the rcv_data and rcv_parity as separate signals,
    // rather than the complete rcv_codeword, because the codeword
    // construction may involve some zero-padded bits that aren't necessary
    // to transmit through the faulty communication channel.
    //
    // The rcv_data is internally zero-padded up to the message size
    // and then concatenated with the rcv_parity to form the received
    // codeword prior to syndrome decoding.
    input  logic                     rcv_valid,
    input  logic [    DataWidth-1:0] rcv_data,
    input  logic [  ParityWidth-1:0] rcv_parity,

    // Decoder output
    output logic                     dec_valid,
    output logic [   InputWidth-1:0] dec_codeword,
    output logic                     dec_error_ce,  // corrected error
    output logic                     dec_error_due,  // detected-but-uncorrectable error
    output logic [  ParityWidth-1:0] dec_error_syndrome,
    output logic [    DataWidth-1:0] dec_data
);

  //------------------------------------------
  // Integration checks
  //------------------------------------------
  `BR_ASSERT_STATIC(data_width_gte_1_a, DataWidth >= 4)
  `BR_ASSERT_STATIC(parity_width_gte_4_a, ParityWidth >= 4)
  `BR_ASSERT_STATIC(parity_width_lte_12_a, ParityWidth <= 12)
  `BR_ASSERT_STATIC(codeword_width_pow_of_2_a, br_math::is_power_of_2(CodewordWidth))
  `BR_ASSERT_STATIC(data_width_fits_in_message_width_a, DataWidth <= MessageWidth)
  `BR_ASSERT_STATIC(right_sized_parity_bits_a, DataWidth > br_ecc::get_max_message_width(ParityWidth - 1))

  //------------------------------------------
  // Implementation
  //------------------------------------------

  //------
  // Optionally register the input signals.
  //------
  logic rcv_valid_d;
  logic [InputWidth-1:0] rcv_codeword_d;

  br_delay_valid #(
      .Width(InputWidth),
      .NumStages(RegisterInputs == 1 ? 1 : 0),
      .EnableAssertFinalNotValid(EnableAssertFinalNotValid)
  ) br_delay_valid_inputs (
      .clk,
      .rst,
      .in_valid(rcv_valid),
      .in({rcv_parity, rcv_data}),
      .out_valid(rcv_valid_d),
      .out(rcv_codeword_d),
      .out_valid_stages(),  // unused
      .out_stages()  // unused
  );

  //------
  // Compute syndrome and set up constant parity check matrix.
  //------
  logic [CodewordWidth-1:0][ParityWidth-1:0] parity_check_matrix;  // H
  logic [ParityWidth-1:0] syndrome;
  logic [CodewordWidth-1:0] cw;  // shorten name for internal readability
  assign `BR_INSERT_TO_MSB(cw, rcv_codeword_d[InputWidth-1 -: ParityWidth])
  if (CodewordWidth > InputWidth) begin : gen_cw_pad_bits
    assign cw[MessageWidth -1 : DataWidth] = '0;
  end
  assign `BR_INSERT_TO_LSB(cw, rcv_codeword_d[DataWidth-1:0])

  // ri lint_check_off EXPR_ID_LIMIT

  if ((CodewordWidth == 8) && (MessageWidth == 4)) begin : gen_8_4
    `BR_ASSERT_STATIC(parity_width_matches_a, ParityWidth == 4)
    assign syndrome[3] = cw[1] ^ cw[2] ^ cw[3] ^ cw[4];
    assign syndrome[2] = cw[0] ^ cw[2] ^ cw[3] ^ cw[5];
    assign syndrome[1] = cw[0] ^ cw[1] ^ cw[3] ^ cw[6];
    assign syndrome[0] = cw[0] ^ cw[1] ^ cw[2] ^ cw[7];
    assign parity_check_matrix[0] = 4'b0111;
    assign parity_check_matrix[1] = 4'b1011;
    assign parity_check_matrix[2] = 4'b1101;
    assign parity_check_matrix[3] = 4'b1110;
    assign parity_check_matrix[4] = 4'b1000;
    assign parity_check_matrix[5] = 4'b0100;
    assign parity_check_matrix[6] = 4'b0010;
    assign parity_check_matrix[7] = 4'b0001;
  end else if ((CodewordWidth == 16) && (MessageWidth == 11)) begin : gen_16_11
    `BR_ASSERT_STATIC(parity_width_matches_a, ParityWidth == 5)
    assign syndrome[4] = cw[0] ^ cw[2] ^ cw[4] ^ cw[5] ^ cw[7] ^ cw[8] ^ cw[10] ^ cw[11];
    assign syndrome[3] = cw[0] ^ cw[2] ^ cw[3] ^ cw[5] ^ cw[6] ^ cw[9] ^ cw[10] ^ cw[12];
    assign syndrome[2] = cw[0] ^ cw[1] ^ cw[3] ^ cw[5] ^ cw[7] ^ cw[8] ^ cw[9] ^ cw[13];
    assign syndrome[1] = cw[0] ^ cw[1] ^ cw[3] ^ cw[4] ^ cw[6] ^ cw[8] ^ cw[10] ^ cw[14];
    assign syndrome[0] = cw[0] ^ cw[1] ^ cw[2] ^ cw[4] ^ cw[6] ^ cw[7] ^ cw[9] ^ cw[15];
    assign parity_check_matrix[0] = 5'b11111;
    assign parity_check_matrix[1] = 5'b00111;
    assign parity_check_matrix[2] = 5'b11001;
    assign parity_check_matrix[3] = 5'b01110;
    assign parity_check_matrix[4] = 5'b10011;
    assign parity_check_matrix[5] = 5'b11100;
    assign parity_check_matrix[6] = 5'b01011;
    assign parity_check_matrix[7] = 5'b10101;
    assign parity_check_matrix[8] = 5'b10110;
    assign parity_check_matrix[9] = 5'b01101;
    assign parity_check_matrix[10] = 5'b11010;
    assign parity_check_matrix[11] = 5'b10000;
    assign parity_check_matrix[12] = 5'b01000;
    assign parity_check_matrix[13] = 5'b00100;
    assign parity_check_matrix[14] = 5'b00010;
    assign parity_check_matrix[15] = 5'b00001;
  end else if ((CodewordWidth == 32) && (MessageWidth == 26)) begin : gen_32_26
    `BR_ASSERT_STATIC(parity_width_matches_a, ParityWidth == 6)
    assign syndrome[5] = cw[1] ^ cw[3] ^ cw[5] ^ cw[6] ^ cw[9] ^ cw[11] ^ cw[12] ^ cw[15] ^ cw[16] ^ cw[18] ^ cw[21] ^ cw[22] ^ cw[23] ^ cw[24] ^ cw[25] ^ cw[26];
    assign syndrome[4] = cw[1] ^ cw[3] ^ cw[4] ^ cw[7] ^ cw[9] ^ cw[10] ^ cw[13] ^ cw[14] ^ cw[17] ^ cw[18] ^ cw[20] ^ cw[22] ^ cw[23] ^ cw[24] ^ cw[25] ^ cw[27];
    assign syndrome[3] = cw[1] ^ cw[2] ^ cw[5] ^ cw[7] ^ cw[8] ^ cw[11] ^ cw[13] ^ cw[14] ^ cw[16] ^ cw[19] ^ cw[20] ^ cw[21] ^ cw[23] ^ cw[24] ^ cw[25] ^ cw[28];
    assign syndrome[2] = cw[0] ^ cw[3] ^ cw[5] ^ cw[7] ^ cw[8] ^ cw[10] ^ cw[12] ^ cw[15] ^ cw[17] ^ cw[19] ^ cw[20] ^ cw[21] ^ cw[22] ^ cw[24] ^ cw[25] ^ cw[29];
    assign syndrome[1] = cw[0] ^ cw[2] ^ cw[4] ^ cw[6] ^ cw[9] ^ cw[11] ^ cw[13] ^ cw[15] ^ cw[17] ^ cw[19] ^ cw[20] ^ cw[21] ^ cw[22] ^ cw[23] ^ cw[25] ^ cw[30];
    assign syndrome[0] = cw[0] ^ cw[2] ^ cw[4] ^ cw[6] ^ cw[8] ^ cw[10] ^ cw[12] ^ cw[14] ^ cw[16] ^ cw[18] ^ cw[20] ^ cw[21] ^ cw[22] ^ cw[23] ^ cw[24] ^ cw[31];
    assign parity_check_matrix[0] = 6'b000111;
    assign parity_check_matrix[1] = 6'b111000;
    assign parity_check_matrix[2] = 6'b001011;
    assign parity_check_matrix[3] = 6'b110100;
    assign parity_check_matrix[4] = 6'b010011;
    assign parity_check_matrix[5] = 6'b101100;
    assign parity_check_matrix[6] = 6'b100011;
    assign parity_check_matrix[7] = 6'b011100;
    assign parity_check_matrix[8] = 6'b001101;
    assign parity_check_matrix[9] = 6'b110010;
    assign parity_check_matrix[10] = 6'b010101;
    assign parity_check_matrix[11] = 6'b101010;
    assign parity_check_matrix[12] = 6'b100101;
    assign parity_check_matrix[13] = 6'b011010;
    assign parity_check_matrix[14] = 6'b011001;
    assign parity_check_matrix[15] = 6'b100110;
    assign parity_check_matrix[16] = 6'b101001;
    assign parity_check_matrix[17] = 6'b010110;
    assign parity_check_matrix[18] = 6'b110001;
    assign parity_check_matrix[19] = 6'b001110;
    assign parity_check_matrix[20] = 6'b011111;
    assign parity_check_matrix[21] = 6'b101111;
    assign parity_check_matrix[22] = 6'b110111;
    assign parity_check_matrix[23] = 6'b111011;
    assign parity_check_matrix[24] = 6'b111101;
    assign parity_check_matrix[25] = 6'b111110;
    assign parity_check_matrix[26] = 6'b100000;
    assign parity_check_matrix[27] = 6'b010000;
    assign parity_check_matrix[28] = 6'b001000;
    assign parity_check_matrix[29] = 6'b000100;
    assign parity_check_matrix[30] = 6'b000010;
    assign parity_check_matrix[31] = 6'b000001;
  end else if ((CodewordWidth == 64) && (MessageWidth == 57)) begin : gen_64_57
    `BR_ASSERT_STATIC(parity_width_matches_a, ParityWidth == 7)
    assign syndrome[6] = cw[0] ^ cw[2] ^ cw[4] ^ cw[6] ^ cw[8] ^ cw[10] ^ cw[12] ^ cw[14] ^ cw[15] ^ cw[17] ^ cw[20] ^ cw[22] ^ cw[24] ^ cw[26] ^ cw[27] ^ cw[30] ^ cw[32] ^ cw[33] ^ cw[35] ^ cw[38] ^ cw[39] ^ cw[42] ^ cw[44] ^ cw[45] ^ cw[47] ^ cw[48] ^ cw[49] ^ cw[50] ^ cw[52] ^ cw[54] ^ cw[56] ^ cw[57];
    assign syndrome[5] = cw[0] ^ cw[2] ^ cw[4] ^ cw[6] ^ cw[8] ^ cw[10] ^ cw[11] ^ cw[13] ^ cw[16] ^ cw[18] ^ cw[20] ^ cw[22] ^ cw[23] ^ cw[26] ^ cw[28] ^ cw[29] ^ cw[31] ^ cw[34] ^ cw[36] ^ cw[38] ^ cw[39] ^ cw[41] ^ cw[43] ^ cw[45] ^ cw[46] ^ cw[49] ^ cw[51] ^ cw[52] ^ cw[54] ^ cw[55] ^ cw[56] ^ cw[58];
    assign syndrome[4] = cw[0] ^ cw[2] ^ cw[4] ^ cw[6] ^ cw[7] ^ cw[9] ^ cw[12] ^ cw[14] ^ cw[16] ^ cw[18] ^ cw[19] ^ cw[22] ^ cw[24] ^ cw[25] ^ cw[28] ^ cw[30] ^ cw[31] ^ cw[34] ^ cw[35] ^ cw[37] ^ cw[40] ^ cw[42] ^ cw[43] ^ cw[45] ^ cw[46] ^ cw[48] ^ cw[50] ^ cw[53] ^ cw[54] ^ cw[55] ^ cw[56] ^ cw[59];
    assign syndrome[3] = cw[0] ^ cw[2] ^ cw[3] ^ cw[5] ^ cw[8] ^ cw[10] ^ cw[12] ^ cw[14] ^ cw[16] ^ cw[18] ^ cw[19] ^ cw[21] ^ cw[23] ^ cw[26] ^ cw[27] ^ cw[30] ^ cw[32] ^ cw[34] ^ cw[36] ^ cw[37] ^ cw[40] ^ cw[41] ^ cw[43] ^ cw[44] ^ cw[47] ^ cw[48] ^ cw[51] ^ cw[52] ^ cw[53] ^ cw[54] ^ cw[56] ^ cw[60];
    assign syndrome[2] = cw[0] ^ cw[1] ^ cw[3] ^ cw[6] ^ cw[7] ^ cw[10] ^ cw[11] ^ cw[14] ^ cw[15] ^ cw[18] ^ cw[20] ^ cw[21] ^ cw[24] ^ cw[25] ^ cw[28] ^ cw[29] ^ cw[32] ^ cw[33] ^ cw[36] ^ cw[38] ^ cw[40] ^ cw[42] ^ cw[43] ^ cw[45] ^ cw[47] ^ cw[48] ^ cw[51] ^ cw[52] ^ cw[53] ^ cw[55] ^ cw[56] ^ cw[61];
    assign syndrome[1] = cw[0] ^ cw[1] ^ cw[3] ^ cw[5] ^ cw[7] ^ cw[9] ^ cw[11] ^ cw[13] ^ cw[15] ^ cw[17] ^ cw[19] ^ cw[22] ^ cw[23] ^ cw[26] ^ cw[27] ^ cw[30] ^ cw[31] ^ cw[34] ^ cw[35] ^ cw[38] ^ cw[39] ^ cw[42] ^ cw[43] ^ cw[45] ^ cw[47] ^ cw[48] ^ cw[51] ^ cw[52] ^ cw[53] ^ cw[54] ^ cw[55] ^ cw[62];
    assign syndrome[0] = cw[0] ^ cw[1] ^ cw[2] ^ cw[5] ^ cw[6] ^ cw[9] ^ cw[10] ^ cw[13] ^ cw[14] ^ cw[17] ^ cw[18] ^ cw[21] ^ cw[22] ^ cw[25] ^ cw[26] ^ cw[29] ^ cw[30] ^ cw[33] ^ cw[34] ^ cw[37] ^ cw[38] ^ cw[41] ^ cw[42] ^ cw[44] ^ cw[46] ^ cw[47] ^ cw[49] ^ cw[50] ^ cw[51] ^ cw[53] ^ cw[55] ^ cw[63];
    assign parity_check_matrix[0] = 7'b1111111;
    assign parity_check_matrix[1] = 7'b0000111;
    assign parity_check_matrix[2] = 7'b1111001;
    assign parity_check_matrix[3] = 7'b0001110;
    assign parity_check_matrix[4] = 7'b1110000;
    assign parity_check_matrix[5] = 7'b0001011;
    assign parity_check_matrix[6] = 7'b1110101;
    assign parity_check_matrix[7] = 7'b0010110;
    assign parity_check_matrix[8] = 7'b1101000;
    assign parity_check_matrix[9] = 7'b0010011;
    assign parity_check_matrix[10] = 7'b1101101;
    assign parity_check_matrix[11] = 7'b0100110;
    assign parity_check_matrix[12] = 7'b1011000;
    assign parity_check_matrix[13] = 7'b0100011;
    assign parity_check_matrix[14] = 7'b1011101;
    assign parity_check_matrix[15] = 7'b1000110;
    assign parity_check_matrix[16] = 7'b0111000;
    assign parity_check_matrix[17] = 7'b1000011;
    assign parity_check_matrix[18] = 7'b0111101;
    assign parity_check_matrix[19] = 7'b0011010;
    assign parity_check_matrix[20] = 7'b1100100;
    assign parity_check_matrix[21] = 7'b0001101;
    assign parity_check_matrix[22] = 7'b1110011;
    assign parity_check_matrix[23] = 7'b0101010;
    assign parity_check_matrix[24] = 7'b1010100;
    assign parity_check_matrix[25] = 7'b0010101;
    assign parity_check_matrix[26] = 7'b1101011;
    assign parity_check_matrix[27] = 7'b1001010;
    assign parity_check_matrix[28] = 7'b0110100;
    assign parity_check_matrix[29] = 7'b0100101;
    assign parity_check_matrix[30] = 7'b1011011;
    assign parity_check_matrix[31] = 7'b0110010;
    assign parity_check_matrix[32] = 7'b1001100;
    assign parity_check_matrix[33] = 7'b1000101;
    assign parity_check_matrix[34] = 7'b0111011;
    assign parity_check_matrix[35] = 7'b1010010;
    assign parity_check_matrix[36] = 7'b0101100;
    assign parity_check_matrix[37] = 7'b0011001;
    assign parity_check_matrix[38] = 7'b1100111;
    assign parity_check_matrix[39] = 7'b1100010;
    assign parity_check_matrix[40] = 7'b0011100;
    assign parity_check_matrix[41] = 7'b0101001;
    assign parity_check_matrix[42] = 7'b1010111;
    assign parity_check_matrix[43] = 7'b0111110;
    assign parity_check_matrix[44] = 7'b1001001;
    assign parity_check_matrix[45] = 7'b1110110;
    assign parity_check_matrix[46] = 7'b0110001;
    assign parity_check_matrix[47] = 7'b1001111;
    assign parity_check_matrix[48] = 7'b1011110;
    assign parity_check_matrix[49] = 7'b1100001;
    assign parity_check_matrix[50] = 7'b1010001;
    assign parity_check_matrix[51] = 7'b0101111;
    assign parity_check_matrix[52] = 7'b1101110;
    assign parity_check_matrix[53] = 7'b0011111;
    assign parity_check_matrix[54] = 7'b1111010;
    assign parity_check_matrix[55] = 7'b0110111;
    assign parity_check_matrix[56] = 7'b1111100;
    assign parity_check_matrix[57] = 7'b1000000;
    assign parity_check_matrix[58] = 7'b0100000;
    assign parity_check_matrix[59] = 7'b0010000;
    assign parity_check_matrix[60] = 7'b0001000;
    assign parity_check_matrix[61] = 7'b0000100;
    assign parity_check_matrix[62] = 7'b0000010;
    assign parity_check_matrix[63] = 7'b0000001;
  end else if ((CodewordWidth == 128) && (MessageWidth == 120)) begin : gen_128_120
    `BR_ASSERT_STATIC(parity_width_matches_a, ParityWidth == 8)
    assign syndrome[7] = cw[1] ^ cw[3] ^ cw[5] ^ cw[7] ^ cw[9] ^ cw[10] ^ cw[13] ^ cw[15] ^ cw[17] ^ cw[19] ^ cw[20] ^ cw[23] ^ cw[25] ^ cw[27] ^ cw[28] ^ cw[31] ^ cw[33] ^ cw[34] ^ cw[37] ^ cw[38] ^ cw[40] ^ cw[43] ^ cw[45] ^ cw[47] ^ cw[49] ^ cw[50] ^ cw[53] ^ cw[55] ^ cw[57] ^ cw[58] ^ cw[61] ^ cw[63] ^ cw[64] ^ cw[67] ^ cw[68] ^ cw[70] ^ cw[73] ^ cw[75] ^ cw[77] ^ cw[78] ^ cw[81] ^ cw[83] ^ cw[84] ^ cw[87] ^ cw[88] ^ cw[90] ^ cw[93] ^ cw[95] ^ cw[96] ^ cw[99] ^ cw[100] ^ cw[102] ^ cw[105] ^ cw[106] ^ cw[108] ^ cw[110] ^ cw[113] ^ cw[114] ^ cw[115] ^ cw[116] ^ cw[117] ^ cw[118] ^ cw[119] ^ cw[120];
    assign syndrome[6] = cw[1] ^ cw[3] ^ cw[5] ^ cw[7] ^ cw[8] ^ cw[11] ^ cw[13] ^ cw[15] ^ cw[17] ^ cw[18] ^ cw[21] ^ cw[23] ^ cw[25] ^ cw[26] ^ cw[29] ^ cw[31] ^ cw[32] ^ cw[35] ^ cw[36] ^ cw[39] ^ cw[40] ^ cw[43] ^ cw[45] ^ cw[47] ^ cw[48] ^ cw[51] ^ cw[53] ^ cw[55] ^ cw[56] ^ cw[59] ^ cw[61] ^ cw[62] ^ cw[65] ^ cw[66] ^ cw[69] ^ cw[70] ^ cw[73] ^ cw[75] ^ cw[76] ^ cw[79] ^ cw[81] ^ cw[82] ^ cw[85] ^ cw[86] ^ cw[89] ^ cw[90] ^ cw[93] ^ cw[94] ^ cw[97] ^ cw[98] ^ cw[101] ^ cw[102] ^ cw[104] ^ cw[107] ^ cw[108] ^ cw[110] ^ cw[112] ^ cw[114] ^ cw[115] ^ cw[116] ^ cw[117] ^ cw[118] ^ cw[119] ^ cw[121];
    assign syndrome[5] = cw[1] ^ cw[3] ^ cw[5] ^ cw[6] ^ cw[9] ^ cw[11] ^ cw[13] ^ cw[15] ^ cw[16] ^ cw[19] ^ cw[21] ^ cw[23] ^ cw[24] ^ cw[27] ^ cw[29] ^ cw[30] ^ cw[33] ^ cw[35] ^ cw[36] ^ cw[38] ^ cw[41] ^ cw[43] ^ cw[45] ^ cw[46] ^ cw[49] ^ cw[51] ^ cw[53] ^ cw[54] ^ cw[57] ^ cw[59] ^ cw[60] ^ cw[63] ^ cw[65] ^ cw[66] ^ cw[68] ^ cw[71] ^ cw[73] ^ cw[74] ^ cw[77] ^ cw[79] ^ cw[80] ^ cw[83] ^ cw[85] ^ cw[86] ^ cw[88] ^ cw[91] ^ cw[92] ^ cw[95] ^ cw[97] ^ cw[98] ^ cw[100] ^ cw[103] ^ cw[104] ^ cw[106] ^ cw[109] ^ cw[110] ^ cw[112] ^ cw[113] ^ cw[115] ^ cw[116] ^ cw[117] ^ cw[118] ^ cw[119] ^ cw[122];
    assign syndrome[4] = cw[1] ^ cw[3] ^ cw[4] ^ cw[7] ^ cw[9] ^ cw[11] ^ cw[13] ^ cw[14] ^ cw[17] ^ cw[19] ^ cw[21] ^ cw[22] ^ cw[25] ^ cw[27] ^ cw[29] ^ cw[30] ^ cw[32] ^ cw[34] ^ cw[37] ^ cw[39] ^ cw[41] ^ cw[43] ^ cw[44] ^ cw[47] ^ cw[49] ^ cw[51] ^ cw[52] ^ cw[55] ^ cw[57] ^ cw[59] ^ cw[60] ^ cw[62] ^ cw[64] ^ cw[67] ^ cw[69] ^ cw[71] ^ cw[72] ^ cw[75] ^ cw[77] ^ cw[79] ^ cw[80] ^ cw[82] ^ cw[84] ^ cw[87] ^ cw[89] ^ cw[91] ^ cw[92] ^ cw[94] ^ cw[96] ^ cw[99] ^ cw[101] ^ cw[103] ^ cw[104] ^ cw[106] ^ cw[108] ^ cw[111] ^ cw[112] ^ cw[113] ^ cw[114] ^ cw[116] ^ cw[117] ^ cw[118] ^ cw[119] ^ cw[123];
    assign syndrome[3] = cw[1] ^ cw[2] ^ cw[5] ^ cw[7] ^ cw[9] ^ cw[11] ^ cw[12] ^ cw[15] ^ cw[17] ^ cw[19] ^ cw[21] ^ cw[22] ^ cw[24] ^ cw[26] ^ cw[28] ^ cw[31] ^ cw[33] ^ cw[35] ^ cw[37] ^ cw[39] ^ cw[41] ^ cw[42] ^ cw[45] ^ cw[47] ^ cw[49] ^ cw[51] ^ cw[52] ^ cw[54] ^ cw[56] ^ cw[58] ^ cw[61] ^ cw[63] ^ cw[65] ^ cw[67] ^ cw[69] ^ cw[71] ^ cw[72] ^ cw[74] ^ cw[76] ^ cw[78] ^ cw[81] ^ cw[83] ^ cw[85] ^ cw[87] ^ cw[89] ^ cw[91] ^ cw[92] ^ cw[94] ^ cw[96] ^ cw[98] ^ cw[100] ^ cw[102] ^ cw[105] ^ cw[107] ^ cw[109] ^ cw[111] ^ cw[112] ^ cw[113] ^ cw[114] ^ cw[115] ^ cw[117] ^ cw[118] ^ cw[119] ^ cw[124];
    assign syndrome[2] = cw[0] ^ cw[3] ^ cw[5] ^ cw[7] ^ cw[9] ^ cw[11] ^ cw[12] ^ cw[14] ^ cw[16] ^ cw[18] ^ cw[20] ^ cw[23] ^ cw[25] ^ cw[27] ^ cw[29] ^ cw[31] ^ cw[33] ^ cw[35] ^ cw[37] ^ cw[39] ^ cw[41] ^ cw[42] ^ cw[44] ^ cw[46] ^ cw[48] ^ cw[50] ^ cw[53] ^ cw[55] ^ cw[57] ^ cw[59] ^ cw[61] ^ cw[63] ^ cw[65] ^ cw[67] ^ cw[69] ^ cw[71] ^ cw[72] ^ cw[74] ^ cw[76] ^ cw[78] ^ cw[80] ^ cw[82] ^ cw[84] ^ cw[86] ^ cw[88] ^ cw[90] ^ cw[93] ^ cw[95] ^ cw[97] ^ cw[99] ^ cw[101] ^ cw[103] ^ cw[105] ^ cw[107] ^ cw[109] ^ cw[111] ^ cw[112] ^ cw[113] ^ cw[114] ^ cw[115] ^ cw[116] ^ cw[118] ^ cw[119] ^ cw[125];
    assign syndrome[1] = cw[0] ^ cw[2] ^ cw[4] ^ cw[6] ^ cw[8] ^ cw[10] ^ cw[13] ^ cw[15] ^ cw[17] ^ cw[19] ^ cw[21] ^ cw[23] ^ cw[25] ^ cw[27] ^ cw[29] ^ cw[31] ^ cw[33] ^ cw[35] ^ cw[37] ^ cw[39] ^ cw[41] ^ cw[42] ^ cw[44] ^ cw[46] ^ cw[48] ^ cw[50] ^ cw[52] ^ cw[54] ^ cw[56] ^ cw[58] ^ cw[60] ^ cw[62] ^ cw[64] ^ cw[66] ^ cw[68] ^ cw[70] ^ cw[73] ^ cw[75] ^ cw[77] ^ cw[79] ^ cw[81] ^ cw[83] ^ cw[85] ^ cw[87] ^ cw[89] ^ cw[91] ^ cw[93] ^ cw[95] ^ cw[97] ^ cw[99] ^ cw[101] ^ cw[103] ^ cw[105] ^ cw[107] ^ cw[109] ^ cw[111] ^ cw[112] ^ cw[113] ^ cw[114] ^ cw[115] ^ cw[116] ^ cw[117] ^ cw[119] ^ cw[126];
    assign syndrome[0] = cw[0] ^ cw[2] ^ cw[4] ^ cw[6] ^ cw[8] ^ cw[10] ^ cw[12] ^ cw[14] ^ cw[16] ^ cw[18] ^ cw[20] ^ cw[22] ^ cw[24] ^ cw[26] ^ cw[28] ^ cw[30] ^ cw[32] ^ cw[34] ^ cw[36] ^ cw[38] ^ cw[40] ^ cw[43] ^ cw[45] ^ cw[47] ^ cw[49] ^ cw[51] ^ cw[53] ^ cw[55] ^ cw[57] ^ cw[59] ^ cw[61] ^ cw[63] ^ cw[65] ^ cw[67] ^ cw[69] ^ cw[71] ^ cw[73] ^ cw[75] ^ cw[77] ^ cw[79] ^ cw[81] ^ cw[83] ^ cw[85] ^ cw[87] ^ cw[89] ^ cw[91] ^ cw[93] ^ cw[95] ^ cw[97] ^ cw[99] ^ cw[101] ^ cw[103] ^ cw[105] ^ cw[107] ^ cw[109] ^ cw[111] ^ cw[112] ^ cw[113] ^ cw[114] ^ cw[115] ^ cw[116] ^ cw[117] ^ cw[118] ^ cw[127];
    assign parity_check_matrix[0] = 8'b00000111;
    assign parity_check_matrix[1] = 8'b11111000;
    assign parity_check_matrix[2] = 8'b00001011;
    assign parity_check_matrix[3] = 8'b11110100;
    assign parity_check_matrix[4] = 8'b00010011;
    assign parity_check_matrix[5] = 8'b11101100;
    assign parity_check_matrix[6] = 8'b00100011;
    assign parity_check_matrix[7] = 8'b11011100;
    assign parity_check_matrix[8] = 8'b01000011;
    assign parity_check_matrix[9] = 8'b10111100;
    assign parity_check_matrix[10] = 8'b10000011;
    assign parity_check_matrix[11] = 8'b01111100;
    assign parity_check_matrix[12] = 8'b00001101;
    assign parity_check_matrix[13] = 8'b11110010;
    assign parity_check_matrix[14] = 8'b00010101;
    assign parity_check_matrix[15] = 8'b11101010;
    assign parity_check_matrix[16] = 8'b00100101;
    assign parity_check_matrix[17] = 8'b11011010;
    assign parity_check_matrix[18] = 8'b01000101;
    assign parity_check_matrix[19] = 8'b10111010;
    assign parity_check_matrix[20] = 8'b10000101;
    assign parity_check_matrix[21] = 8'b01111010;
    assign parity_check_matrix[22] = 8'b00011001;
    assign parity_check_matrix[23] = 8'b11100110;
    assign parity_check_matrix[24] = 8'b00101001;
    assign parity_check_matrix[25] = 8'b11010110;
    assign parity_check_matrix[26] = 8'b01001001;
    assign parity_check_matrix[27] = 8'b10110110;
    assign parity_check_matrix[28] = 8'b10001001;
    assign parity_check_matrix[29] = 8'b01110110;
    assign parity_check_matrix[30] = 8'b00110001;
    assign parity_check_matrix[31] = 8'b11001110;
    assign parity_check_matrix[32] = 8'b01010001;
    assign parity_check_matrix[33] = 8'b10101110;
    assign parity_check_matrix[34] = 8'b10010001;
    assign parity_check_matrix[35] = 8'b01101110;
    assign parity_check_matrix[36] = 8'b01100001;
    assign parity_check_matrix[37] = 8'b10011110;
    assign parity_check_matrix[38] = 8'b10100001;
    assign parity_check_matrix[39] = 8'b01011110;
    assign parity_check_matrix[40] = 8'b11000001;
    assign parity_check_matrix[41] = 8'b00111110;
    assign parity_check_matrix[42] = 8'b00001110;
    assign parity_check_matrix[43] = 8'b11110001;
    assign parity_check_matrix[44] = 8'b00010110;
    assign parity_check_matrix[45] = 8'b11101001;
    assign parity_check_matrix[46] = 8'b00100110;
    assign parity_check_matrix[47] = 8'b11011001;
    assign parity_check_matrix[48] = 8'b01000110;
    assign parity_check_matrix[49] = 8'b10111001;
    assign parity_check_matrix[50] = 8'b10000110;
    assign parity_check_matrix[51] = 8'b01111001;
    assign parity_check_matrix[52] = 8'b00011010;
    assign parity_check_matrix[53] = 8'b11100101;
    assign parity_check_matrix[54] = 8'b00101010;
    assign parity_check_matrix[55] = 8'b11010101;
    assign parity_check_matrix[56] = 8'b01001010;
    assign parity_check_matrix[57] = 8'b10110101;
    assign parity_check_matrix[58] = 8'b10001010;
    assign parity_check_matrix[59] = 8'b01110101;
    assign parity_check_matrix[60] = 8'b00110010;
    assign parity_check_matrix[61] = 8'b11001101;
    assign parity_check_matrix[62] = 8'b01010010;
    assign parity_check_matrix[63] = 8'b10101101;
    assign parity_check_matrix[64] = 8'b10010010;
    assign parity_check_matrix[65] = 8'b01101101;
    assign parity_check_matrix[66] = 8'b01100010;
    assign parity_check_matrix[67] = 8'b10011101;
    assign parity_check_matrix[68] = 8'b10100010;
    assign parity_check_matrix[69] = 8'b01011101;
    assign parity_check_matrix[70] = 8'b11000010;
    assign parity_check_matrix[71] = 8'b00111101;
    assign parity_check_matrix[72] = 8'b00011100;
    assign parity_check_matrix[73] = 8'b11100011;
    assign parity_check_matrix[74] = 8'b00101100;
    assign parity_check_matrix[75] = 8'b11010011;
    assign parity_check_matrix[76] = 8'b01001100;
    assign parity_check_matrix[77] = 8'b10110011;
    assign parity_check_matrix[78] = 8'b10001100;
    assign parity_check_matrix[79] = 8'b01110011;
    assign parity_check_matrix[80] = 8'b00110100;
    assign parity_check_matrix[81] = 8'b11001011;
    assign parity_check_matrix[82] = 8'b01010100;
    assign parity_check_matrix[83] = 8'b10101011;
    assign parity_check_matrix[84] = 8'b10010100;
    assign parity_check_matrix[85] = 8'b01101011;
    assign parity_check_matrix[86] = 8'b01100100;
    assign parity_check_matrix[87] = 8'b10011011;
    assign parity_check_matrix[88] = 8'b10100100;
    assign parity_check_matrix[89] = 8'b01011011;
    assign parity_check_matrix[90] = 8'b11000100;
    assign parity_check_matrix[91] = 8'b00111011;
    assign parity_check_matrix[92] = 8'b00111000;
    assign parity_check_matrix[93] = 8'b11000111;
    assign parity_check_matrix[94] = 8'b01011000;
    assign parity_check_matrix[95] = 8'b10100111;
    assign parity_check_matrix[96] = 8'b10011000;
    assign parity_check_matrix[97] = 8'b01100111;
    assign parity_check_matrix[98] = 8'b01101000;
    assign parity_check_matrix[99] = 8'b10010111;
    assign parity_check_matrix[100] = 8'b10101000;
    assign parity_check_matrix[101] = 8'b01010111;
    assign parity_check_matrix[102] = 8'b11001000;
    assign parity_check_matrix[103] = 8'b00110111;
    assign parity_check_matrix[104] = 8'b01110000;
    assign parity_check_matrix[105] = 8'b10001111;
    assign parity_check_matrix[106] = 8'b10110000;
    assign parity_check_matrix[107] = 8'b01001111;
    assign parity_check_matrix[108] = 8'b11010000;
    assign parity_check_matrix[109] = 8'b00101111;
    assign parity_check_matrix[110] = 8'b11100000;
    assign parity_check_matrix[111] = 8'b00011111;
    assign parity_check_matrix[112] = 8'b01111111;
    assign parity_check_matrix[113] = 8'b10111111;
    assign parity_check_matrix[114] = 8'b11011111;
    assign parity_check_matrix[115] = 8'b11101111;
    assign parity_check_matrix[116] = 8'b11110111;
    assign parity_check_matrix[117] = 8'b11111011;
    assign parity_check_matrix[118] = 8'b11111101;
    assign parity_check_matrix[119] = 8'b11111110;
    assign parity_check_matrix[120] = 8'b10000000;
    assign parity_check_matrix[121] = 8'b01000000;
    assign parity_check_matrix[122] = 8'b00100000;
    assign parity_check_matrix[123] = 8'b00010000;
    assign parity_check_matrix[124] = 8'b00001000;
    assign parity_check_matrix[125] = 8'b00000100;
    assign parity_check_matrix[126] = 8'b00000010;
    assign parity_check_matrix[127] = 8'b00000001;
  end else if ((CodewordWidth == 256) && (MessageWidth == 247)) begin : gen_256_247
    `BR_ASSERT_STATIC(parity_width_matches_a, ParityWidth == 9)
    assign syndrome[8] = cw[0] ^ cw[2] ^ cw[4] ^ cw[6] ^ cw[8] ^ cw[10] ^ cw[12] ^ cw[14] ^ cw[16] ^ cw[18] ^ cw[20] ^ cw[22] ^ cw[23] ^ cw[25] ^ cw[28] ^ cw[30] ^ cw[32] ^ cw[34] ^ cw[36] ^ cw[38] ^ cw[40] ^ cw[42] ^ cw[43] ^ cw[46] ^ cw[48] ^ cw[49] ^ cw[52] ^ cw[54] ^ cw[56] ^ cw[58] ^ cw[59] ^ cw[62] ^ cw[64] ^ cw[66] ^ cw[68] ^ cw[69] ^ cw[71] ^ cw[74] ^ cw[76] ^ cw[78] ^ cw[79] ^ cw[82] ^ cw[83] ^ cw[85] ^ cw[88] ^ cw[90] ^ cw[92] ^ cw[94] ^ cw[96] ^ cw[97] ^ cw[100] ^ cw[102] ^ cw[103] ^ cw[105] ^ cw[108] ^ cw[109] ^ cw[112] ^ cw[115] ^ cw[117] ^ cw[119] ^ cw[120] ^ cw[124] ^ cw[126] ^ cw[129] ^ cw[130] ^ cw[132] ^ cw[135] ^ cw[137] ^ cw[139] ^ cw[143] ^ cw[144] ^ cw[147] ^ cw[148] ^ cw[152] ^ cw[153] ^ cw[155] ^ cw[158] ^ cw[159] ^ cw[161] ^ cw[162] ^ cw[166] ^ cw[168] ^ cw[170] ^ cw[171] ^ cw[173] ^ cw[175] ^ cw[177] ^ cw[178] ^ cw[180] ^ cw[181] ^ cw[183] ^ cw[185] ^ cw[187] ^ cw[188] ^ cw[190] ^ cw[193] ^ cw[194] ^ cw[195] ^ cw[198] ^ cw[200] ^ cw[201] ^ cw[203] ^ cw[205] ^ cw[206] ^ cw[209] ^ cw[211] ^ cw[212] ^ cw[214] ^ cw[215] ^ cw[218] ^ cw[220] ^ cw[221] ^ cw[223] ^ cw[225] ^ cw[227] ^ cw[228] ^ cw[230] ^ cw[232] ^ cw[234] ^ cw[236] ^ cw[237] ^ cw[239] ^ cw[240] ^ cw[242] ^ cw[243] ^ cw[245] ^ cw[246] ^ cw[247];
    assign syndrome[7] = cw[0] ^ cw[2] ^ cw[4] ^ cw[6] ^ cw[8] ^ cw[10] ^ cw[12] ^ cw[14] ^ cw[16] ^ cw[18] ^ cw[19] ^ cw[21] ^ cw[24] ^ cw[26] ^ cw[28] ^ cw[30] ^ cw[32] ^ cw[34] ^ cw[36] ^ cw[38] ^ cw[39] ^ cw[42] ^ cw[44] ^ cw[45] ^ cw[48] ^ cw[50] ^ cw[52] ^ cw[54] ^ cw[55] ^ cw[58] ^ cw[60] ^ cw[62] ^ cw[64] ^ cw[65] ^ cw[67] ^ cw[70] ^ cw[72] ^ cw[74] ^ cw[75] ^ cw[78] ^ cw[80] ^ cw[81] ^ cw[83] ^ cw[86] ^ cw[88] ^ cw[90] ^ cw[92] ^ cw[93] ^ cw[96] ^ cw[98] ^ cw[99] ^ cw[101] ^ cw[104] ^ cw[106] ^ cw[108] ^ cw[109] ^ cw[112] ^ cw[113] ^ cw[117] ^ cw[119] ^ cw[121] ^ cw[123] ^ cw[126] ^ cw[128] ^ cw[131] ^ cw[133] ^ cw[134] ^ cw[138] ^ cw[140] ^ cw[141] ^ cw[144] ^ cw[146] ^ cw[148] ^ cw[150] ^ cw[153] ^ cw[154] ^ cw[156] ^ cw[159] ^ cw[161] ^ cw[163] ^ cw[164] ^ cw[168] ^ cw[170] ^ cw[171] ^ cw[173] ^ cw[175] ^ cw[177] ^ cw[178] ^ cw[179] ^ cw[181] ^ cw[182] ^ cw[184] ^ cw[186] ^ cw[189] ^ cw[191] ^ cw[193] ^ cw[194] ^ cw[196] ^ cw[198] ^ cw[199] ^ cw[201] ^ cw[202] ^ cw[204] ^ cw[207] ^ cw[208] ^ cw[210] ^ cw[212] ^ cw[214] ^ cw[216] ^ cw[218] ^ cw[219] ^ cw[222] ^ cw[224] ^ cw[226] ^ cw[227] ^ cw[229] ^ cw[230] ^ cw[233] ^ cw[234] ^ cw[236] ^ cw[238] ^ cw[239] ^ cw[241] ^ cw[242] ^ cw[244] ^ cw[245] ^ cw[246] ^ cw[248];
    assign syndrome[6] = cw[0] ^ cw[2] ^ cw[4] ^ cw[6] ^ cw[8] ^ cw[10] ^ cw[12] ^ cw[14] ^ cw[15] ^ cw[17] ^ cw[20] ^ cw[22] ^ cw[24] ^ cw[26] ^ cw[28] ^ cw[30] ^ cw[32] ^ cw[34] ^ cw[35] ^ cw[38] ^ cw[40] ^ cw[41] ^ cw[44] ^ cw[46] ^ cw[48] ^ cw[50] ^ cw[51] ^ cw[54] ^ cw[56] ^ cw[58] ^ cw[60] ^ cw[61] ^ cw[63] ^ cw[66] ^ cw[68] ^ cw[70] ^ cw[72] ^ cw[74] ^ cw[75] ^ cw[77] ^ cw[79] ^ cw[82] ^ cw[84] ^ cw[86] ^ cw[88] ^ cw[89] ^ cw[92] ^ cw[94] ^ cw[95] ^ cw[98] ^ cw[100] ^ cw[101] ^ cw[104] ^ cw[105] ^ cw[108] ^ cw[110] ^ cw[111] ^ cw[114] ^ cw[116] ^ cw[119] ^ cw[122] ^ cw[124] ^ cw[125] ^ cw[127] ^ cw[131] ^ cw[133] ^ cw[135] ^ cw[138] ^ cw[140] ^ cw[141] ^ cw[143] ^ cw[146] ^ cw[149] ^ cw[150] ^ cw[152] ^ cw[154] ^ cw[157] ^ cw[158] ^ cw[161] ^ cw[162] ^ cw[165] ^ cw[167] ^ cw[170] ^ cw[171] ^ cw[172] ^ cw[174] ^ cw[176] ^ cw[178] ^ cw[180] ^ cw[181] ^ cw[183] ^ cw[185] ^ cw[187] ^ cw[189] ^ cw[191] ^ cw[192] ^ cw[194] ^ cw[196] ^ cw[197] ^ cw[200] ^ cw[201] ^ cw[203] ^ cw[204] ^ cw[207] ^ cw[208] ^ cw[211] ^ cw[212] ^ cw[213] ^ cw[215] ^ cw[217] ^ cw[220] ^ cw[222] ^ cw[223] ^ cw[225] ^ cw[226] ^ cw[229] ^ cw[231] ^ cw[232] ^ cw[234] ^ cw[235] ^ cw[238] ^ cw[239] ^ cw[240] ^ cw[241] ^ cw[243] ^ cw[244] ^ cw[245] ^ cw[249];
    assign syndrome[5] = cw[0] ^ cw[2] ^ cw[4] ^ cw[6] ^ cw[8] ^ cw[10] ^ cw[11] ^ cw[13] ^ cw[16] ^ cw[18] ^ cw[20] ^ cw[22] ^ cw[24] ^ cw[26] ^ cw[28] ^ cw[30] ^ cw[31] ^ cw[34] ^ cw[36] ^ cw[37] ^ cw[40] ^ cw[42] ^ cw[44] ^ cw[46] ^ cw[47] ^ cw[50] ^ cw[52] ^ cw[54] ^ cw[56] ^ cw[57] ^ cw[60] ^ cw[62] ^ cw[63] ^ cw[66] ^ cw[67] ^ cw[70] ^ cw[71] ^ cw[73] ^ cw[76] ^ cw[78] ^ cw[80] ^ cw[82] ^ cw[84] ^ cw[86] ^ cw[88] ^ cw[89] ^ cw[91] ^ cw[93] ^ cw[96] ^ cw[97] ^ cw[100] ^ cw[102] ^ cw[104] ^ cw[106] ^ cw[107] ^ cw[110] ^ cw[112] ^ cw[114] ^ cw[116] ^ cw[118] ^ cw[121] ^ cw[123] ^ cw[126] ^ cw[127] ^ cw[130] ^ cw[133] ^ cw[134] ^ cw[137] ^ cw[139] ^ cw[142] ^ cw[145] ^ cw[147] ^ cw[150] ^ cw[151] ^ cw[155] ^ cw[157] ^ cw[158] ^ cw[159] ^ cw[160] ^ cw[162] ^ cw[166] ^ cw[168] ^ cw[169] ^ cw[171] ^ cw[172] ^ cw[175] ^ cw[176] ^ cw[178] ^ cw[180] ^ cw[181] ^ cw[182] ^ cw[185] ^ cw[186] ^ cw[189] ^ cw[191] ^ cw[192] ^ cw[194] ^ cw[196] ^ cw[197] ^ cw[199] ^ cw[201] ^ cw[202] ^ cw[205] ^ cw[206] ^ cw[209] ^ cw[210] ^ cw[211] ^ cw[213] ^ cw[216] ^ cw[217] ^ cw[219] ^ cw[221] ^ cw[224] ^ cw[226] ^ cw[227] ^ cw[228] ^ cw[231] ^ cw[232] ^ cw[233] ^ cw[235] ^ cw[237] ^ cw[238] ^ cw[240] ^ cw[242] ^ cw[243] ^ cw[244] ^ cw[246] ^ cw[250];
    assign syndrome[4] = cw[0] ^ cw[2] ^ cw[4] ^ cw[6] ^ cw[7] ^ cw[9] ^ cw[12] ^ cw[14] ^ cw[16] ^ cw[18] ^ cw[20] ^ cw[22] ^ cw[24] ^ cw[26] ^ cw[27] ^ cw[30] ^ cw[32] ^ cw[33] ^ cw[36] ^ cw[38] ^ cw[40] ^ cw[42] ^ cw[44] ^ cw[46] ^ cw[47] ^ cw[50] ^ cw[51] ^ cw[53] ^ cw[55] ^ cw[58] ^ cw[59] ^ cw[62] ^ cw[64] ^ cw[66] ^ cw[68] ^ cw[70] ^ cw[72] ^ cw[73] ^ cw[76] ^ cw[77] ^ cw[80] ^ cw[81] ^ cw[84] ^ cw[85] ^ cw[87] ^ cw[90] ^ cw[92] ^ cw[94] ^ cw[96] ^ cw[98] ^ cw[100] ^ cw[102] ^ cw[104] ^ cw[106] ^ cw[107] ^ cw[110] ^ cw[111] ^ cw[113] ^ cw[116] ^ cw[118] ^ cw[120] ^ cw[123] ^ cw[125] ^ cw[128] ^ cw[129] ^ cw[132] ^ cw[136] ^ cw[137] ^ cw[140] ^ cw[142] ^ cw[145] ^ cw[147] ^ cw[149] ^ cw[152] ^ cw[153] ^ cw[154] ^ cw[158] ^ cw[160] ^ cw[163] ^ cw[164] ^ cw[165] ^ cw[167] ^ cw[169] ^ cw[171] ^ cw[173] ^ cw[174] ^ cw[176] ^ cw[178] ^ cw[179] ^ cw[181] ^ cw[183] ^ cw[184] ^ cw[186] ^ cw[188] ^ cw[190] ^ cw[192] ^ cw[193] ^ cw[195] ^ cw[196] ^ cw[199] ^ cw[200] ^ cw[203] ^ cw[205] ^ cw[206] ^ cw[208] ^ cw[211] ^ cw[212] ^ cw[213] ^ cw[214] ^ cw[216] ^ cw[220] ^ cw[222] ^ cw[224] ^ cw[225] ^ cw[227] ^ cw[228] ^ cw[229] ^ cw[230] ^ cw[231] ^ cw[233] ^ cw[235] ^ cw[236] ^ cw[237] ^ cw[241] ^ cw[244] ^ cw[245] ^ cw[246] ^ cw[251];
    assign syndrome[3] = cw[0] ^ cw[2] ^ cw[3] ^ cw[5] ^ cw[8] ^ cw[10] ^ cw[12] ^ cw[14] ^ cw[16] ^ cw[18] ^ cw[20] ^ cw[22] ^ cw[24] ^ cw[26] ^ cw[27] ^ cw[29] ^ cw[31] ^ cw[34] ^ cw[35] ^ cw[38] ^ cw[39] ^ cw[42] ^ cw[43] ^ cw[46] ^ cw[48] ^ cw[50] ^ cw[52] ^ cw[53] ^ cw[56] ^ cw[57] ^ cw[60] ^ cw[61] ^ cw[64] ^ cw[65] ^ cw[68] ^ cw[69] ^ cw[72] ^ cw[74] ^ cw[76] ^ cw[78] ^ cw[80] ^ cw[82] ^ cw[84] ^ cw[86] ^ cw[87] ^ cw[90] ^ cw[91] ^ cw[94] ^ cw[95] ^ cw[98] ^ cw[99] ^ cw[102] ^ cw[103] ^ cw[106] ^ cw[108] ^ cw[110] ^ cw[112] ^ cw[114] ^ cw[115] ^ cw[118] ^ cw[121] ^ cw[122] ^ cw[125] ^ cw[128] ^ cw[130] ^ cw[132] ^ cw[135] ^ cw[136] ^ cw[138] ^ cw[142] ^ cw[144] ^ cw[146] ^ cw[149] ^ cw[151] ^ cw[156] ^ cw[157] ^ cw[158] ^ cw[160] ^ cw[164] ^ cw[165] ^ cw[166] ^ cw[168] ^ cw[169] ^ cw[171] ^ cw[173] ^ cw[174] ^ cw[176] ^ cw[177] ^ cw[179] ^ cw[181] ^ cw[183] ^ cw[184] ^ cw[186] ^ cw[187] ^ cw[188] ^ cw[190] ^ cw[191] ^ cw[194] ^ cw[195] ^ cw[197] ^ cw[198] ^ cw[202] ^ cw[204] ^ cw[206] ^ cw[207] ^ cw[208] ^ cw[209] ^ cw[210] ^ cw[212] ^ cw[215] ^ cw[217] ^ cw[218] ^ cw[219] ^ cw[221] ^ cw[223] ^ cw[225] ^ cw[226] ^ cw[230] ^ cw[232] ^ cw[233] ^ cw[235] ^ cw[237] ^ cw[239] ^ cw[241] ^ cw[243] ^ cw[244] ^ cw[246] ^ cw[252];
    assign syndrome[2] = cw[0] ^ cw[1] ^ cw[3] ^ cw[6] ^ cw[7] ^ cw[10] ^ cw[11] ^ cw[14] ^ cw[15] ^ cw[18] ^ cw[19] ^ cw[22] ^ cw[23] ^ cw[26] ^ cw[28] ^ cw[29] ^ cw[32] ^ cw[33] ^ cw[36] ^ cw[37] ^ cw[40] ^ cw[41] ^ cw[44] ^ cw[45] ^ cw[48] ^ cw[49] ^ cw[52] ^ cw[54] ^ cw[56] ^ cw[58] ^ cw[60] ^ cw[62] ^ cw[64] ^ cw[66] ^ cw[68] ^ cw[70] ^ cw[72] ^ cw[74] ^ cw[76] ^ cw[78] ^ cw[80] ^ cw[82] ^ cw[84] ^ cw[86] ^ cw[87] ^ cw[90] ^ cw[91] ^ cw[94] ^ cw[95] ^ cw[98] ^ cw[99] ^ cw[102] ^ cw[103] ^ cw[106] ^ cw[107] ^ cw[110] ^ cw[111] ^ cw[113] ^ cw[115] ^ cw[117] ^ cw[120] ^ cw[122] ^ cw[124] ^ cw[127] ^ cw[129] ^ cw[131] ^ cw[134] ^ cw[136] ^ cw[139] ^ cw[141] ^ cw[143] ^ cw[145] ^ cw[148] ^ cw[151] ^ cw[155] ^ cw[156] ^ cw[158] ^ cw[160] ^ cw[163] ^ cw[165] ^ cw[166] ^ cw[167] ^ cw[169] ^ cw[170] ^ cw[172] ^ cw[174] ^ cw[175] ^ cw[178] ^ cw[179] ^ cw[181] ^ cw[182] ^ cw[184] ^ cw[185] ^ cw[189] ^ cw[190] ^ cw[192] ^ cw[194] ^ cw[195] ^ cw[197] ^ cw[198] ^ cw[199] ^ cw[202] ^ cw[203] ^ cw[204] ^ cw[205] ^ cw[207] ^ cw[212] ^ cw[214] ^ cw[215] ^ cw[217] ^ cw[218] ^ cw[219] ^ cw[220] ^ cw[221] ^ cw[222] ^ cw[223] ^ cw[224] ^ cw[228] ^ cw[229] ^ cw[231] ^ cw[234] ^ cw[236] ^ cw[238] ^ cw[240] ^ cw[242] ^ cw[244] ^ cw[246] ^ cw[253];
    assign syndrome[1] = cw[0] ^ cw[1] ^ cw[3] ^ cw[5] ^ cw[7] ^ cw[9] ^ cw[11] ^ cw[13] ^ cw[15] ^ cw[17] ^ cw[19] ^ cw[21] ^ cw[23] ^ cw[25] ^ cw[27] ^ cw[30] ^ cw[31] ^ cw[34] ^ cw[35] ^ cw[38] ^ cw[39] ^ cw[42] ^ cw[43] ^ cw[46] ^ cw[47] ^ cw[50] ^ cw[51] ^ cw[54] ^ cw[55] ^ cw[58] ^ cw[59] ^ cw[62] ^ cw[63] ^ cw[66] ^ cw[67] ^ cw[70] ^ cw[71] ^ cw[74] ^ cw[75] ^ cw[78] ^ cw[79] ^ cw[82] ^ cw[83] ^ cw[86] ^ cw[88] ^ cw[90] ^ cw[92] ^ cw[94] ^ cw[96] ^ cw[98] ^ cw[100] ^ cw[102] ^ cw[104] ^ cw[106] ^ cw[108] ^ cw[110] ^ cw[112] ^ cw[115] ^ cw[117] ^ cw[119] ^ cw[122] ^ cw[124] ^ cw[126] ^ cw[129] ^ cw[131] ^ cw[133] ^ cw[136] ^ cw[138] ^ cw[140] ^ cw[142] ^ cw[145] ^ cw[147] ^ cw[149] ^ cw[151] ^ cw[155] ^ cw[156] ^ cw[157] ^ cw[158] ^ cw[163] ^ cw[164] ^ cw[166] ^ cw[167] ^ cw[169] ^ cw[171] ^ cw[172] ^ cw[174] ^ cw[176] ^ cw[177] ^ cw[178] ^ cw[180] ^ cw[182] ^ cw[184] ^ cw[186] ^ cw[187] ^ cw[188] ^ cw[190] ^ cw[192] ^ cw[193] ^ cw[194] ^ cw[197] ^ cw[199] ^ cw[200] ^ cw[202] ^ cw[204] ^ cw[206] ^ cw[208] ^ cw[209] ^ cw[210] ^ cw[212] ^ cw[213] ^ cw[215] ^ cw[216] ^ cw[218] ^ cw[220] ^ cw[222] ^ cw[225] ^ cw[226] ^ cw[228] ^ cw[230] ^ cw[232] ^ cw[234] ^ cw[236] ^ cw[238] ^ cw[240] ^ cw[242] ^ cw[244] ^ cw[246] ^ cw[254];
    assign syndrome[0] = cw[0] ^ cw[1] ^ cw[2] ^ cw[5] ^ cw[6] ^ cw[9] ^ cw[10] ^ cw[13] ^ cw[14] ^ cw[17] ^ cw[18] ^ cw[21] ^ cw[22] ^ cw[25] ^ cw[26] ^ cw[29] ^ cw[30] ^ cw[33] ^ cw[34] ^ cw[37] ^ cw[38] ^ cw[41] ^ cw[42] ^ cw[45] ^ cw[46] ^ cw[49] ^ cw[50] ^ cw[53] ^ cw[54] ^ cw[57] ^ cw[58] ^ cw[61] ^ cw[62] ^ cw[65] ^ cw[66] ^ cw[69] ^ cw[70] ^ cw[73] ^ cw[74] ^ cw[77] ^ cw[78] ^ cw[81] ^ cw[82] ^ cw[85] ^ cw[86] ^ cw[89] ^ cw[90] ^ cw[93] ^ cw[94] ^ cw[97] ^ cw[98] ^ cw[101] ^ cw[102] ^ cw[105] ^ cw[106] ^ cw[109] ^ cw[110] ^ cw[115] ^ cw[117] ^ cw[119] ^ cw[122] ^ cw[124] ^ cw[126] ^ cw[129] ^ cw[131] ^ cw[133] ^ cw[136] ^ cw[138] ^ cw[140] ^ cw[142] ^ cw[145] ^ cw[147] ^ cw[149] ^ cw[151] ^ cw[155] ^ cw[156] ^ cw[157] ^ cw[160] ^ cw[163] ^ cw[164] ^ cw[165] ^ cw[167] ^ cw[168] ^ cw[170] ^ cw[172] ^ cw[173] ^ cw[175] ^ cw[177] ^ cw[179] ^ cw[180] ^ cw[182] ^ cw[183] ^ cw[185] ^ cw[187] ^ cw[188] ^ cw[189] ^ cw[191] ^ cw[193] ^ cw[195] ^ cw[196] ^ cw[198] ^ cw[200] ^ cw[201] ^ cw[203] ^ cw[205] ^ cw[207] ^ cw[209] ^ cw[210] ^ cw[211] ^ cw[213] ^ cw[214] ^ cw[216] ^ cw[217] ^ cw[219] ^ cw[221] ^ cw[223] ^ cw[224] ^ cw[227] ^ cw[229] ^ cw[231] ^ cw[233] ^ cw[235] ^ cw[237] ^ cw[239] ^ cw[241] ^ cw[243] ^ cw[245] ^ cw[255];
    assign parity_check_matrix[0] = 9'b111111111;
    assign parity_check_matrix[1] = 9'b000000111;
    assign parity_check_matrix[2] = 9'b111111001;
    assign parity_check_matrix[3] = 9'b000001110;
    assign parity_check_matrix[4] = 9'b111110000;
    assign parity_check_matrix[5] = 9'b000001011;
    assign parity_check_matrix[6] = 9'b111110101;
    assign parity_check_matrix[7] = 9'b000010110;
    assign parity_check_matrix[8] = 9'b111101000;
    assign parity_check_matrix[9] = 9'b000010011;
    assign parity_check_matrix[10] = 9'b111101101;
    assign parity_check_matrix[11] = 9'b000100110;
    assign parity_check_matrix[12] = 9'b111011000;
    assign parity_check_matrix[13] = 9'b000100011;
    assign parity_check_matrix[14] = 9'b111011101;
    assign parity_check_matrix[15] = 9'b001000110;
    assign parity_check_matrix[16] = 9'b110111000;
    assign parity_check_matrix[17] = 9'b001000011;
    assign parity_check_matrix[18] = 9'b110111101;
    assign parity_check_matrix[19] = 9'b010000110;
    assign parity_check_matrix[20] = 9'b101111000;
    assign parity_check_matrix[21] = 9'b010000011;
    assign parity_check_matrix[22] = 9'b101111101;
    assign parity_check_matrix[23] = 9'b100000110;
    assign parity_check_matrix[24] = 9'b011111000;
    assign parity_check_matrix[25] = 9'b100000011;
    assign parity_check_matrix[26] = 9'b011111101;
    assign parity_check_matrix[27] = 9'b000011010;
    assign parity_check_matrix[28] = 9'b111100100;
    assign parity_check_matrix[29] = 9'b000001101;
    assign parity_check_matrix[30] = 9'b111110011;
    assign parity_check_matrix[31] = 9'b000101010;
    assign parity_check_matrix[32] = 9'b111010100;
    assign parity_check_matrix[33] = 9'b000010101;
    assign parity_check_matrix[34] = 9'b111101011;
    assign parity_check_matrix[35] = 9'b001001010;
    assign parity_check_matrix[36] = 9'b110110100;
    assign parity_check_matrix[37] = 9'b000100101;
    assign parity_check_matrix[38] = 9'b111011011;
    assign parity_check_matrix[39] = 9'b010001010;
    assign parity_check_matrix[40] = 9'b101110100;
    assign parity_check_matrix[41] = 9'b001000101;
    assign parity_check_matrix[42] = 9'b110111011;
    assign parity_check_matrix[43] = 9'b100001010;
    assign parity_check_matrix[44] = 9'b011110100;
    assign parity_check_matrix[45] = 9'b010000101;
    assign parity_check_matrix[46] = 9'b101111011;
    assign parity_check_matrix[47] = 9'b000110010;
    assign parity_check_matrix[48] = 9'b111001100;
    assign parity_check_matrix[49] = 9'b100000101;
    assign parity_check_matrix[50] = 9'b011111011;
    assign parity_check_matrix[51] = 9'b001010010;
    assign parity_check_matrix[52] = 9'b110101100;
    assign parity_check_matrix[53] = 9'b000011001;
    assign parity_check_matrix[54] = 9'b111100111;
    assign parity_check_matrix[55] = 9'b010010010;
    assign parity_check_matrix[56] = 9'b101101100;
    assign parity_check_matrix[57] = 9'b000101001;
    assign parity_check_matrix[58] = 9'b111010111;
    assign parity_check_matrix[59] = 9'b100010010;
    assign parity_check_matrix[60] = 9'b011101100;
    assign parity_check_matrix[61] = 9'b001001001;
    assign parity_check_matrix[62] = 9'b110110111;
    assign parity_check_matrix[63] = 9'b001100010;
    assign parity_check_matrix[64] = 9'b110011100;
    assign parity_check_matrix[65] = 9'b010001001;
    assign parity_check_matrix[66] = 9'b101110111;
    assign parity_check_matrix[67] = 9'b010100010;
    assign parity_check_matrix[68] = 9'b101011100;
    assign parity_check_matrix[69] = 9'b100001001;
    assign parity_check_matrix[70] = 9'b011110111;
    assign parity_check_matrix[71] = 9'b100100010;
    assign parity_check_matrix[72] = 9'b011011100;
    assign parity_check_matrix[73] = 9'b000110001;
    assign parity_check_matrix[74] = 9'b111001111;
    assign parity_check_matrix[75] = 9'b011000010;
    assign parity_check_matrix[76] = 9'b100111100;
    assign parity_check_matrix[77] = 9'b001010001;
    assign parity_check_matrix[78] = 9'b110101111;
    assign parity_check_matrix[79] = 9'b101000010;
    assign parity_check_matrix[80] = 9'b010111100;
    assign parity_check_matrix[81] = 9'b010010001;
    assign parity_check_matrix[82] = 9'b101101111;
    assign parity_check_matrix[83] = 9'b110000010;
    assign parity_check_matrix[84] = 9'b001111100;
    assign parity_check_matrix[85] = 9'b100010001;
    assign parity_check_matrix[86] = 9'b011101111;
    assign parity_check_matrix[87] = 9'b000011100;
    assign parity_check_matrix[88] = 9'b111100010;
    assign parity_check_matrix[89] = 9'b001100001;
    assign parity_check_matrix[90] = 9'b110011111;
    assign parity_check_matrix[91] = 9'b000101100;
    assign parity_check_matrix[92] = 9'b111010010;
    assign parity_check_matrix[93] = 9'b010100001;
    assign parity_check_matrix[94] = 9'b101011111;
    assign parity_check_matrix[95] = 9'b001001100;
    assign parity_check_matrix[96] = 9'b110110010;
    assign parity_check_matrix[97] = 9'b100100001;
    assign parity_check_matrix[98] = 9'b011011111;
    assign parity_check_matrix[99] = 9'b010001100;
    assign parity_check_matrix[100] = 9'b101110010;
    assign parity_check_matrix[101] = 9'b011000001;
    assign parity_check_matrix[102] = 9'b100111111;
    assign parity_check_matrix[103] = 9'b100001100;
    assign parity_check_matrix[104] = 9'b011110010;
    assign parity_check_matrix[105] = 9'b101000001;
    assign parity_check_matrix[106] = 9'b010111111;
    assign parity_check_matrix[107] = 9'b000110100;
    assign parity_check_matrix[108] = 9'b111001010;
    assign parity_check_matrix[109] = 9'b110000001;
    assign parity_check_matrix[110] = 9'b001111111;
    assign parity_check_matrix[111] = 9'b001010100;
    assign parity_check_matrix[112] = 9'b110101010;
    assign parity_check_matrix[113] = 9'b010010100;
    assign parity_check_matrix[114] = 9'b001101000;
    assign parity_check_matrix[115] = 9'b100001111;
    assign parity_check_matrix[116] = 9'b001110000;
    assign parity_check_matrix[117] = 9'b110000111;
    assign parity_check_matrix[118] = 9'b000111000;
    assign parity_check_matrix[119] = 9'b111000011;
    assign parity_check_matrix[120] = 9'b100010100;
    assign parity_check_matrix[121] = 9'b010101000;
    assign parity_check_matrix[122] = 9'b001001111;
    assign parity_check_matrix[123] = 9'b010110000;
    assign parity_check_matrix[124] = 9'b101000111;
    assign parity_check_matrix[125] = 9'b001011000;
    assign parity_check_matrix[126] = 9'b110100011;
    assign parity_check_matrix[127] = 9'b001100100;
    assign parity_check_matrix[128] = 9'b010011000;
    assign parity_check_matrix[129] = 9'b100010111;
    assign parity_check_matrix[130] = 9'b100101000;
    assign parity_check_matrix[131] = 9'b011000111;
    assign parity_check_matrix[132] = 9'b100011000;
    assign parity_check_matrix[133] = 9'b011100011;
    assign parity_check_matrix[134] = 9'b010100100;
    assign parity_check_matrix[135] = 9'b101001000;
    assign parity_check_matrix[136] = 9'b000011111;
    assign parity_check_matrix[137] = 9'b100110000;
    assign parity_check_matrix[138] = 9'b011001011;
    assign parity_check_matrix[139] = 9'b100100100;
    assign parity_check_matrix[140] = 9'b011010011;
    assign parity_check_matrix[141] = 9'b011000100;
    assign parity_check_matrix[142] = 9'b000111011;
    assign parity_check_matrix[143] = 9'b101000100;
    assign parity_check_matrix[144] = 9'b110001000;
    assign parity_check_matrix[145] = 9'b000110111;
    assign parity_check_matrix[146] = 9'b011001000;
    assign parity_check_matrix[147] = 9'b100110011;
    assign parity_check_matrix[148] = 9'b110000100;
    assign parity_check_matrix[149] = 9'b001011011;
    assign parity_check_matrix[150] = 9'b011100000;
    assign parity_check_matrix[151] = 9'b000101111;
    assign parity_check_matrix[152] = 9'b101010000;
    assign parity_check_matrix[153] = 9'b110010000;
    assign parity_check_matrix[154] = 9'b011010000;
    assign parity_check_matrix[155] = 9'b100100111;
    assign parity_check_matrix[156] = 9'b010001111;
    assign parity_check_matrix[157] = 9'b001101011;
    assign parity_check_matrix[158] = 9'b101111110;
    assign parity_check_matrix[159] = 9'b110100000;
    assign parity_check_matrix[160] = 9'b000111101;
    assign parity_check_matrix[161] = 9'b111000000;
    assign parity_check_matrix[162] = 9'b101100000;
    assign parity_check_matrix[163] = 9'b010010111;
    assign parity_check_matrix[164] = 9'b010011011;
    assign parity_check_matrix[165] = 9'b001011101;
    assign parity_check_matrix[166] = 9'b100101110;
    assign parity_check_matrix[167] = 9'b001010111;
    assign parity_check_matrix[168] = 9'b110101001;
    assign parity_check_matrix[169] = 9'b000111110;
    assign parity_check_matrix[170] = 9'b111000101;
    assign parity_check_matrix[171] = 9'b111111010;
    assign parity_check_matrix[172] = 9'b001100111;
    assign parity_check_matrix[173] = 9'b110011001;
    assign parity_check_matrix[174] = 9'b001011110;
    assign parity_check_matrix[175] = 9'b110100101;
    assign parity_check_matrix[176] = 9'b001111010;
    assign parity_check_matrix[177] = 9'b110001011;
    assign parity_check_matrix[178] = 9'b111110110;
    assign parity_check_matrix[179] = 9'b010011101;
    assign parity_check_matrix[180] = 9'b101100011;
    assign parity_check_matrix[181] = 9'b111111100;
    assign parity_check_matrix[182] = 9'b010100111;
    assign parity_check_matrix[183] = 9'b101011001;
    assign parity_check_matrix[184] = 9'b010011110;
    assign parity_check_matrix[185] = 9'b101100101;
    assign parity_check_matrix[186] = 9'b010111010;
    assign parity_check_matrix[187] = 9'b101001011;
    assign parity_check_matrix[188] = 9'b100011011;
    assign parity_check_matrix[189] = 9'b011100101;
    assign parity_check_matrix[190] = 9'b100011110;
    assign parity_check_matrix[191] = 9'b011101001;
    assign parity_check_matrix[192] = 9'b001110110;
    assign parity_check_matrix[193] = 9'b110010011;
    assign parity_check_matrix[194] = 9'b111101110;
    assign parity_check_matrix[195] = 9'b100011101;
    assign parity_check_matrix[196] = 9'b011110001;
    assign parity_check_matrix[197] = 9'b001101110;
    assign parity_check_matrix[198] = 9'b110001101;
    assign parity_check_matrix[199] = 9'b010110110;
    assign parity_check_matrix[200] = 9'b101010011;
    assign parity_check_matrix[201] = 9'b111100001;
    assign parity_check_matrix[202] = 9'b010101110;
    assign parity_check_matrix[203] = 9'b101010101;
    assign parity_check_matrix[204] = 9'b011001110;
    assign parity_check_matrix[205] = 9'b100110101;
    assign parity_check_matrix[206] = 9'b100111010;
    assign parity_check_matrix[207] = 9'b011001101;
    assign parity_check_matrix[208] = 9'b011011010;
    assign parity_check_matrix[209] = 9'b100101011;
    assign parity_check_matrix[210] = 9'b010101011;
    assign parity_check_matrix[211] = 9'b101110001;
    assign parity_check_matrix[212] = 9'b111011110;
    assign parity_check_matrix[213] = 9'b001110011;
    assign parity_check_matrix[214] = 9'b110010101;
    assign parity_check_matrix[215] = 9'b101001110;
    assign parity_check_matrix[216] = 9'b010110011;
    assign parity_check_matrix[217] = 9'b001101101;
    assign parity_check_matrix[218] = 9'b110001110;
    assign parity_check_matrix[219] = 9'b010101101;
    assign parity_check_matrix[220] = 9'b101010110;
    assign parity_check_matrix[221] = 9'b100101101;
    assign parity_check_matrix[222] = 9'b011010110;
    assign parity_check_matrix[223] = 9'b101001101;
    assign parity_check_matrix[224] = 9'b010110101;
    assign parity_check_matrix[225] = 9'b101011010;
    assign parity_check_matrix[226] = 9'b011101010;
    assign parity_check_matrix[227] = 9'b110110001;
    assign parity_check_matrix[228] = 9'b100110110;
    assign parity_check_matrix[229] = 9'b011010101;
    assign parity_check_matrix[230] = 9'b110011010;
    assign parity_check_matrix[231] = 9'b001110101;
    assign parity_check_matrix[232] = 9'b101101010;
    assign parity_check_matrix[233] = 9'b010111001;
    assign parity_check_matrix[234] = 9'b111000110;
    assign parity_check_matrix[235] = 9'b001111001;
    assign parity_check_matrix[236] = 9'b110010110;
    assign parity_check_matrix[237] = 9'b100111001;
    assign parity_check_matrix[238] = 9'b011100110;
    assign parity_check_matrix[239] = 9'b111001001;
    assign parity_check_matrix[240] = 9'b101100110;
    assign parity_check_matrix[241] = 9'b011011001;
    assign parity_check_matrix[242] = 9'b110100110;
    assign parity_check_matrix[243] = 9'b101101001;
    assign parity_check_matrix[244] = 9'b011111110;
    assign parity_check_matrix[245] = 9'b111010001;
    assign parity_check_matrix[246] = 9'b110111110;
    assign parity_check_matrix[247] = 9'b100000000;
    assign parity_check_matrix[248] = 9'b010000000;
    assign parity_check_matrix[249] = 9'b001000000;
    assign parity_check_matrix[250] = 9'b000100000;
    assign parity_check_matrix[251] = 9'b000010000;
    assign parity_check_matrix[252] = 9'b000001000;
    assign parity_check_matrix[253] = 9'b000000100;
    assign parity_check_matrix[254] = 9'b000000010;
    assign parity_check_matrix[255] = 9'b000000001;
  end else if ((CodewordWidth == 512) && (MessageWidth == 502)) begin : gen_512_502
    `BR_ASSERT_STATIC(parity_width_matches_a, ParityWidth == 10)
    assign syndrome[9] = cw[1] ^ cw[3] ^ cw[5] ^ cw[7] ^ cw[9] ^ cw[11] ^ cw[13] ^ cw[14] ^ cw[17] ^ cw[19] ^ cw[21] ^ cw[23] ^ cw[25] ^ cw[27] ^ cw[28] ^ cw[31] ^ cw[33] ^ cw[35] ^ cw[37] ^ cw[39] ^ cw[40] ^ cw[43] ^ cw[45] ^ cw[47] ^ cw[49] ^ cw[50] ^ cw[53] ^ cw[55] ^ cw[57] ^ cw[58] ^ cw[61] ^ cw[63] ^ cw[64] ^ cw[67] ^ cw[68] ^ cw[70] ^ cw[73] ^ cw[75] ^ cw[77] ^ cw[79] ^ cw[81] ^ cw[83] ^ cw[84] ^ cw[87] ^ cw[89] ^ cw[91] ^ cw[93] ^ cw[95] ^ cw[96] ^ cw[99] ^ cw[101] ^ cw[103] ^ cw[105] ^ cw[106] ^ cw[109] ^ cw[111] ^ cw[113] ^ cw[114] ^ cw[117] ^ cw[119] ^ cw[120] ^ cw[123] ^ cw[124] ^ cw[126] ^ cw[129] ^ cw[131] ^ cw[133] ^ cw[135] ^ cw[137] ^ cw[138] ^ cw[141] ^ cw[143] ^ cw[145] ^ cw[147] ^ cw[148] ^ cw[151] ^ cw[153] ^ cw[155] ^ cw[156] ^ cw[159] ^ cw[161] ^ cw[162] ^ cw[165] ^ cw[166] ^ cw[168] ^ cw[171] ^ cw[173] ^ cw[175] ^ cw[177] ^ cw[178] ^ cw[181] ^ cw[183] ^ cw[185] ^ cw[186] ^ cw[189] ^ cw[191] ^ cw[192] ^ cw[195] ^ cw[196] ^ cw[198] ^ cw[201] ^ cw[203] ^ cw[205] ^ cw[206] ^ cw[209] ^ cw[211] ^ cw[212] ^ cw[215] ^ cw[216] ^ cw[218] ^ cw[221] ^ cw[223] ^ cw[224] ^ cw[227] ^ cw[228] ^ cw[230] ^ cw[233] ^ cw[234] ^ cw[236] ^ cw[238] ^ cw[241] ^ cw[243] ^ cw[245] ^ cw[247] ^ cw[249] ^ cw[250] ^ cw[253] ^ cw[255] ^ cw[257] ^ cw[259] ^ cw[260] ^ cw[263] ^ cw[265] ^ cw[267] ^ cw[268] ^ cw[271] ^ cw[273] ^ cw[274] ^ cw[277] ^ cw[278] ^ cw[280] ^ cw[283] ^ cw[285] ^ cw[287] ^ cw[289] ^ cw[290] ^ cw[293] ^ cw[295] ^ cw[297] ^ cw[298] ^ cw[301] ^ cw[303] ^ cw[304] ^ cw[307] ^ cw[308] ^ cw[310] ^ cw[313] ^ cw[315] ^ cw[317] ^ cw[318] ^ cw[321] ^ cw[323] ^ cw[324] ^ cw[327] ^ cw[328] ^ cw[330] ^ cw[333] ^ cw[335] ^ cw[336] ^ cw[339] ^ cw[340] ^ cw[342] ^ cw[345] ^ cw[346] ^ cw[348] ^ cw[350] ^ cw[353] ^ cw[355] ^ cw[357] ^ cw[359] ^ cw[360] ^ cw[363] ^ cw[365] ^ cw[367] ^ cw[368] ^ cw[371] ^ cw[373] ^ cw[374] ^ cw[377] ^ cw[378] ^ cw[380] ^ cw[383] ^ cw[385] ^ cw[387] ^ cw[388] ^ cw[391] ^ cw[393] ^ cw[394] ^ cw[397] ^ cw[398] ^ cw[400] ^ cw[403] ^ cw[405] ^ cw[406] ^ cw[409] ^ cw[410] ^ cw[412] ^ cw[415] ^ cw[416] ^ cw[418] ^ cw[420] ^ cw[423] ^ cw[425] ^ cw[427] ^ cw[428] ^ cw[431] ^ cw[433] ^ cw[434] ^ cw[437] ^ cw[438] ^ cw[440] ^ cw[443] ^ cw[445] ^ cw[446] ^ cw[449] ^ cw[450] ^ cw[452] ^ cw[455] ^ cw[456] ^ cw[458] ^ cw[460] ^ cw[463] ^ cw[465] ^ cw[466] ^ cw[469] ^ cw[470] ^ cw[472] ^ cw[475] ^ cw[476] ^ cw[478] ^ cw[480] ^ cw[483] ^ cw[484] ^ cw[486] ^ cw[488] ^ cw[490] ^ cw[493] ^ cw[494] ^ cw[495] ^ cw[496] ^ cw[497] ^ cw[498] ^ cw[499] ^ cw[500] ^ cw[501] ^ cw[502];
    assign syndrome[8] = cw[1] ^ cw[3] ^ cw[5] ^ cw[7] ^ cw[9] ^ cw[11] ^ cw[12] ^ cw[15] ^ cw[17] ^ cw[19] ^ cw[21] ^ cw[23] ^ cw[25] ^ cw[26] ^ cw[29] ^ cw[31] ^ cw[33] ^ cw[35] ^ cw[37] ^ cw[38] ^ cw[41] ^ cw[43] ^ cw[45] ^ cw[47] ^ cw[48] ^ cw[51] ^ cw[53] ^ cw[55] ^ cw[56] ^ cw[59] ^ cw[61] ^ cw[62] ^ cw[65] ^ cw[66] ^ cw[69] ^ cw[70] ^ cw[73] ^ cw[75] ^ cw[77] ^ cw[79] ^ cw[81] ^ cw[82] ^ cw[85] ^ cw[87] ^ cw[89] ^ cw[91] ^ cw[93] ^ cw[94] ^ cw[97] ^ cw[99] ^ cw[101] ^ cw[103] ^ cw[104] ^ cw[107] ^ cw[109] ^ cw[111] ^ cw[112] ^ cw[115] ^ cw[117] ^ cw[118] ^ cw[121] ^ cw[122] ^ cw[125] ^ cw[126] ^ cw[129] ^ cw[131] ^ cw[133] ^ cw[135] ^ cw[136] ^ cw[139] ^ cw[141] ^ cw[143] ^ cw[145] ^ cw[146] ^ cw[149] ^ cw[151] ^ cw[153] ^ cw[154] ^ cw[157] ^ cw[159] ^ cw[160] ^ cw[163] ^ cw[164] ^ cw[167] ^ cw[168] ^ cw[171] ^ cw[173] ^ cw[175] ^ cw[176] ^ cw[179] ^ cw[181] ^ cw[183] ^ cw[184] ^ cw[187] ^ cw[189] ^ cw[190] ^ cw[193] ^ cw[194] ^ cw[197] ^ cw[198] ^ cw[201] ^ cw[203] ^ cw[204] ^ cw[207] ^ cw[209] ^ cw[210] ^ cw[213] ^ cw[214] ^ cw[217] ^ cw[218] ^ cw[221] ^ cw[222] ^ cw[225] ^ cw[226] ^ cw[229] ^ cw[230] ^ cw[232] ^ cw[235] ^ cw[236] ^ cw[238] ^ cw[241] ^ cw[243] ^ cw[245] ^ cw[247] ^ cw[248] ^ cw[251] ^ cw[253] ^ cw[255] ^ cw[257] ^ cw[258] ^ cw[261] ^ cw[263] ^ cw[265] ^ cw[266] ^ cw[269] ^ cw[271] ^ cw[272] ^ cw[275] ^ cw[276] ^ cw[279] ^ cw[280] ^ cw[283] ^ cw[285] ^ cw[287] ^ cw[288] ^ cw[291] ^ cw[293] ^ cw[295] ^ cw[296] ^ cw[299] ^ cw[301] ^ cw[302] ^ cw[305] ^ cw[306] ^ cw[309] ^ cw[310] ^ cw[313] ^ cw[315] ^ cw[316] ^ cw[319] ^ cw[321] ^ cw[322] ^ cw[325] ^ cw[326] ^ cw[329] ^ cw[330] ^ cw[333] ^ cw[334] ^ cw[337] ^ cw[338] ^ cw[341] ^ cw[342] ^ cw[344] ^ cw[347] ^ cw[348] ^ cw[350] ^ cw[353] ^ cw[355] ^ cw[357] ^ cw[358] ^ cw[361] ^ cw[363] ^ cw[365] ^ cw[366] ^ cw[369] ^ cw[371] ^ cw[372] ^ cw[375] ^ cw[376] ^ cw[379] ^ cw[380] ^ cw[383] ^ cw[385] ^ cw[386] ^ cw[389] ^ cw[391] ^ cw[392] ^ cw[395] ^ cw[396] ^ cw[399] ^ cw[400] ^ cw[403] ^ cw[404] ^ cw[407] ^ cw[408] ^ cw[411] ^ cw[412] ^ cw[414] ^ cw[417] ^ cw[418] ^ cw[420] ^ cw[423] ^ cw[425] ^ cw[426] ^ cw[429] ^ cw[431] ^ cw[432] ^ cw[435] ^ cw[436] ^ cw[439] ^ cw[440] ^ cw[443] ^ cw[444] ^ cw[447] ^ cw[448] ^ cw[451] ^ cw[452] ^ cw[454] ^ cw[457] ^ cw[458] ^ cw[460] ^ cw[463] ^ cw[464] ^ cw[467] ^ cw[468] ^ cw[471] ^ cw[472] ^ cw[474] ^ cw[477] ^ cw[478] ^ cw[480] ^ cw[482] ^ cw[485] ^ cw[486] ^ cw[488] ^ cw[490] ^ cw[492] ^ cw[494] ^ cw[495] ^ cw[496] ^ cw[497] ^ cw[498] ^ cw[499] ^ cw[500] ^ cw[501] ^ cw[503];
    assign syndrome[7] = cw[1] ^ cw[3] ^ cw[5] ^ cw[7] ^ cw[9] ^ cw[10] ^ cw[13] ^ cw[15] ^ cw[17] ^ cw[19] ^ cw[21] ^ cw[23] ^ cw[24] ^ cw[27] ^ cw[29] ^ cw[31] ^ cw[33] ^ cw[35] ^ cw[36] ^ cw[39] ^ cw[41] ^ cw[43] ^ cw[45] ^ cw[46] ^ cw[49] ^ cw[51] ^ cw[53] ^ cw[54] ^ cw[57] ^ cw[59] ^ cw[60] ^ cw[63] ^ cw[65] ^ cw[66] ^ cw[68] ^ cw[71] ^ cw[73] ^ cw[75] ^ cw[77] ^ cw[79] ^ cw[80] ^ cw[83] ^ cw[85] ^ cw[87] ^ cw[89] ^ cw[91] ^ cw[92] ^ cw[95] ^ cw[97] ^ cw[99] ^ cw[101] ^ cw[102] ^ cw[105] ^ cw[107] ^ cw[109] ^ cw[110] ^ cw[113] ^ cw[115] ^ cw[116] ^ cw[119] ^ cw[121] ^ cw[122] ^ cw[124] ^ cw[127] ^ cw[129] ^ cw[131] ^ cw[133] ^ cw[134] ^ cw[137] ^ cw[139] ^ cw[141] ^ cw[143] ^ cw[144] ^ cw[147] ^ cw[149] ^ cw[151] ^ cw[152] ^ cw[155] ^ cw[157] ^ cw[158] ^ cw[161] ^ cw[163] ^ cw[164] ^ cw[166] ^ cw[169] ^ cw[171] ^ cw[173] ^ cw[174] ^ cw[177] ^ cw[179] ^ cw[181] ^ cw[182] ^ cw[185] ^ cw[187] ^ cw[188] ^ cw[191] ^ cw[193] ^ cw[194] ^ cw[196] ^ cw[199] ^ cw[201] ^ cw[202] ^ cw[205] ^ cw[207] ^ cw[208] ^ cw[211] ^ cw[213] ^ cw[214] ^ cw[216] ^ cw[219] ^ cw[220] ^ cw[223] ^ cw[225] ^ cw[226] ^ cw[228] ^ cw[231] ^ cw[232] ^ cw[234] ^ cw[237] ^ cw[238] ^ cw[241] ^ cw[243] ^ cw[245] ^ cw[246] ^ cw[249] ^ cw[251] ^ cw[253] ^ cw[255] ^ cw[256] ^ cw[259] ^ cw[261] ^ cw[263] ^ cw[264] ^ cw[267] ^ cw[269] ^ cw[270] ^ cw[273] ^ cw[275] ^ cw[276] ^ cw[278] ^ cw[281] ^ cw[283] ^ cw[285] ^ cw[286] ^ cw[289] ^ cw[291] ^ cw[293] ^ cw[294] ^ cw[297] ^ cw[299] ^ cw[300] ^ cw[303] ^ cw[305] ^ cw[306] ^ cw[308] ^ cw[311] ^ cw[313] ^ cw[314] ^ cw[317] ^ cw[319] ^ cw[320] ^ cw[323] ^ cw[325] ^ cw[326] ^ cw[328] ^ cw[331] ^ cw[332] ^ cw[335] ^ cw[337] ^ cw[338] ^ cw[340] ^ cw[343] ^ cw[344] ^ cw[346] ^ cw[349] ^ cw[350] ^ cw[353] ^ cw[355] ^ cw[356] ^ cw[359] ^ cw[361] ^ cw[363] ^ cw[364] ^ cw[367] ^ cw[369] ^ cw[370] ^ cw[373] ^ cw[375] ^ cw[376] ^ cw[378] ^ cw[381] ^ cw[383] ^ cw[384] ^ cw[387] ^ cw[389] ^ cw[390] ^ cw[393] ^ cw[395] ^ cw[396] ^ cw[398] ^ cw[401] ^ cw[402] ^ cw[405] ^ cw[407] ^ cw[408] ^ cw[410] ^ cw[413] ^ cw[414] ^ cw[416] ^ cw[419] ^ cw[420] ^ cw[423] ^ cw[424] ^ cw[427] ^ cw[429] ^ cw[430] ^ cw[433] ^ cw[435] ^ cw[436] ^ cw[438] ^ cw[441] ^ cw[442] ^ cw[445] ^ cw[447] ^ cw[448] ^ cw[450] ^ cw[453] ^ cw[454] ^ cw[456] ^ cw[459] ^ cw[460] ^ cw[462] ^ cw[465] ^ cw[467] ^ cw[468] ^ cw[470] ^ cw[473] ^ cw[474] ^ cw[476] ^ cw[479] ^ cw[480] ^ cw[482] ^ cw[484] ^ cw[487] ^ cw[488] ^ cw[490] ^ cw[492] ^ cw[493] ^ cw[495] ^ cw[496] ^ cw[497] ^ cw[498] ^ cw[499] ^ cw[500] ^ cw[501] ^ cw[504];
    assign syndrome[6] = cw[1] ^ cw[3] ^ cw[5] ^ cw[7] ^ cw[8] ^ cw[11] ^ cw[13] ^ cw[15] ^ cw[17] ^ cw[19] ^ cw[21] ^ cw[22] ^ cw[25] ^ cw[27] ^ cw[29] ^ cw[31] ^ cw[33] ^ cw[34] ^ cw[37] ^ cw[39] ^ cw[41] ^ cw[43] ^ cw[44] ^ cw[47] ^ cw[49] ^ cw[51] ^ cw[52] ^ cw[55] ^ cw[57] ^ cw[59] ^ cw[60] ^ cw[62] ^ cw[64] ^ cw[67] ^ cw[69] ^ cw[71] ^ cw[73] ^ cw[75] ^ cw[77] ^ cw[78] ^ cw[81] ^ cw[83] ^ cw[85] ^ cw[87] ^ cw[89] ^ cw[90] ^ cw[93] ^ cw[95] ^ cw[97] ^ cw[99] ^ cw[100] ^ cw[103] ^ cw[105] ^ cw[107] ^ cw[108] ^ cw[111] ^ cw[113] ^ cw[115] ^ cw[116] ^ cw[118] ^ cw[120] ^ cw[123] ^ cw[125] ^ cw[127] ^ cw[129] ^ cw[131] ^ cw[132] ^ cw[135] ^ cw[137] ^ cw[139] ^ cw[141] ^ cw[142] ^ cw[145] ^ cw[147] ^ cw[149] ^ cw[150] ^ cw[153] ^ cw[155] ^ cw[157] ^ cw[158] ^ cw[160] ^ cw[162] ^ cw[165] ^ cw[167] ^ cw[169] ^ cw[171] ^ cw[172] ^ cw[175] ^ cw[177] ^ cw[179] ^ cw[180] ^ cw[183] ^ cw[185] ^ cw[187] ^ cw[188] ^ cw[190] ^ cw[192] ^ cw[195] ^ cw[197] ^ cw[199] ^ cw[200] ^ cw[203] ^ cw[205] ^ cw[207] ^ cw[208] ^ cw[210] ^ cw[212] ^ cw[215] ^ cw[217] ^ cw[219] ^ cw[220] ^ cw[222] ^ cw[224] ^ cw[227] ^ cw[229] ^ cw[231] ^ cw[232] ^ cw[234] ^ cw[236] ^ cw[239] ^ cw[241] ^ cw[243] ^ cw[244] ^ cw[247] ^ cw[249] ^ cw[251] ^ cw[253] ^ cw[254] ^ cw[257] ^ cw[259] ^ cw[261] ^ cw[262] ^ cw[265] ^ cw[267] ^ cw[269] ^ cw[270] ^ cw[272] ^ cw[274] ^ cw[277] ^ cw[279] ^ cw[281] ^ cw[283] ^ cw[284] ^ cw[287] ^ cw[289] ^ cw[291] ^ cw[292] ^ cw[295] ^ cw[297] ^ cw[299] ^ cw[300] ^ cw[302] ^ cw[304] ^ cw[307] ^ cw[309] ^ cw[311] ^ cw[312] ^ cw[315] ^ cw[317] ^ cw[319] ^ cw[320] ^ cw[322] ^ cw[324] ^ cw[327] ^ cw[329] ^ cw[331] ^ cw[332] ^ cw[334] ^ cw[336] ^ cw[339] ^ cw[341] ^ cw[343] ^ cw[344] ^ cw[346] ^ cw[348] ^ cw[351] ^ cw[353] ^ cw[354] ^ cw[357] ^ cw[359] ^ cw[361] ^ cw[362] ^ cw[365] ^ cw[367] ^ cw[369] ^ cw[370] ^ cw[372] ^ cw[374] ^ cw[377] ^ cw[379] ^ cw[381] ^ cw[382] ^ cw[385] ^ cw[387] ^ cw[389] ^ cw[390] ^ cw[392] ^ cw[394] ^ cw[397] ^ cw[399] ^ cw[401] ^ cw[402] ^ cw[404] ^ cw[406] ^ cw[409] ^ cw[411] ^ cw[413] ^ cw[414] ^ cw[416] ^ cw[418] ^ cw[421] ^ cw[422] ^ cw[425] ^ cw[427] ^ cw[429] ^ cw[430] ^ cw[432] ^ cw[434] ^ cw[437] ^ cw[439] ^ cw[441] ^ cw[442] ^ cw[444] ^ cw[446] ^ cw[449] ^ cw[451] ^ cw[453] ^ cw[454] ^ cw[456] ^ cw[458] ^ cw[461] ^ cw[462] ^ cw[464] ^ cw[466] ^ cw[469] ^ cw[471] ^ cw[473] ^ cw[474] ^ cw[476] ^ cw[478] ^ cw[481] ^ cw[482] ^ cw[484] ^ cw[486] ^ cw[489] ^ cw[490] ^ cw[492] ^ cw[493] ^ cw[494] ^ cw[496] ^ cw[497] ^ cw[498] ^ cw[499] ^ cw[500] ^ cw[501] ^ cw[505];
    assign syndrome[5] = cw[1] ^ cw[3] ^ cw[5] ^ cw[6] ^ cw[9] ^ cw[11] ^ cw[13] ^ cw[15] ^ cw[17] ^ cw[19] ^ cw[20] ^ cw[23] ^ cw[25] ^ cw[27] ^ cw[29] ^ cw[31] ^ cw[32] ^ cw[35] ^ cw[37] ^ cw[39] ^ cw[41] ^ cw[42] ^ cw[45] ^ cw[47] ^ cw[49] ^ cw[51] ^ cw[52] ^ cw[54] ^ cw[56] ^ cw[58] ^ cw[61] ^ cw[63] ^ cw[65] ^ cw[67] ^ cw[69] ^ cw[71] ^ cw[73] ^ cw[75] ^ cw[76] ^ cw[79] ^ cw[81] ^ cw[83] ^ cw[85] ^ cw[87] ^ cw[88] ^ cw[91] ^ cw[93] ^ cw[95] ^ cw[97] ^ cw[98] ^ cw[101] ^ cw[103] ^ cw[105] ^ cw[107] ^ cw[108] ^ cw[110] ^ cw[112] ^ cw[114] ^ cw[117] ^ cw[119] ^ cw[121] ^ cw[123] ^ cw[125] ^ cw[127] ^ cw[129] ^ cw[130] ^ cw[133] ^ cw[135] ^ cw[137] ^ cw[139] ^ cw[140] ^ cw[143] ^ cw[145] ^ cw[147] ^ cw[149] ^ cw[150] ^ cw[152] ^ cw[154] ^ cw[156] ^ cw[159] ^ cw[161] ^ cw[163] ^ cw[165] ^ cw[167] ^ cw[169] ^ cw[170] ^ cw[173] ^ cw[175] ^ cw[177] ^ cw[179] ^ cw[180] ^ cw[182] ^ cw[184] ^ cw[186] ^ cw[189] ^ cw[191] ^ cw[193] ^ cw[195] ^ cw[197] ^ cw[199] ^ cw[200] ^ cw[202] ^ cw[204] ^ cw[206] ^ cw[209] ^ cw[211] ^ cw[213] ^ cw[215] ^ cw[217] ^ cw[219] ^ cw[220] ^ cw[222] ^ cw[224] ^ cw[226] ^ cw[228] ^ cw[230] ^ cw[233] ^ cw[235] ^ cw[237] ^ cw[239] ^ cw[241] ^ cw[242] ^ cw[245] ^ cw[247] ^ cw[249] ^ cw[251] ^ cw[252] ^ cw[255] ^ cw[257] ^ cw[259] ^ cw[261] ^ cw[262] ^ cw[264] ^ cw[266] ^ cw[268] ^ cw[271] ^ cw[273] ^ cw[275] ^ cw[277] ^ cw[279] ^ cw[281] ^ cw[282] ^ cw[285] ^ cw[287] ^ cw[289] ^ cw[291] ^ cw[292] ^ cw[294] ^ cw[296] ^ cw[298] ^ cw[301] ^ cw[303] ^ cw[305] ^ cw[307] ^ cw[309] ^ cw[311] ^ cw[312] ^ cw[314] ^ cw[316] ^ cw[318] ^ cw[321] ^ cw[323] ^ cw[325] ^ cw[327] ^ cw[329] ^ cw[331] ^ cw[332] ^ cw[334] ^ cw[336] ^ cw[338] ^ cw[340] ^ cw[342] ^ cw[345] ^ cw[347] ^ cw[349] ^ cw[351] ^ cw[352] ^ cw[355] ^ cw[357] ^ cw[359] ^ cw[361] ^ cw[362] ^ cw[364] ^ cw[366] ^ cw[368] ^ cw[371] ^ cw[373] ^ cw[375] ^ cw[377] ^ cw[379] ^ cw[381] ^ cw[382] ^ cw[384] ^ cw[386] ^ cw[388] ^ cw[391] ^ cw[393] ^ cw[395] ^ cw[397] ^ cw[399] ^ cw[401] ^ cw[402] ^ cw[404] ^ cw[406] ^ cw[408] ^ cw[410] ^ cw[412] ^ cw[415] ^ cw[417] ^ cw[419] ^ cw[421] ^ cw[422] ^ cw[424] ^ cw[426] ^ cw[428] ^ cw[431] ^ cw[433] ^ cw[435] ^ cw[437] ^ cw[439] ^ cw[441] ^ cw[442] ^ cw[444] ^ cw[446] ^ cw[448] ^ cw[450] ^ cw[452] ^ cw[455] ^ cw[457] ^ cw[459] ^ cw[461] ^ cw[462] ^ cw[464] ^ cw[466] ^ cw[468] ^ cw[470] ^ cw[472] ^ cw[475] ^ cw[477] ^ cw[479] ^ cw[481] ^ cw[482] ^ cw[484] ^ cw[486] ^ cw[488] ^ cw[491] ^ cw[492] ^ cw[493] ^ cw[494] ^ cw[495] ^ cw[497] ^ cw[498] ^ cw[499] ^ cw[500] ^ cw[501] ^ cw[506];
    assign syndrome[4] = cw[1] ^ cw[3] ^ cw[4] ^ cw[7] ^ cw[9] ^ cw[11] ^ cw[13] ^ cw[15] ^ cw[17] ^ cw[18] ^ cw[21] ^ cw[23] ^ cw[25] ^ cw[27] ^ cw[29] ^ cw[30] ^ cw[33] ^ cw[35] ^ cw[37] ^ cw[39] ^ cw[41] ^ cw[42] ^ cw[44] ^ cw[46] ^ cw[48] ^ cw[50] ^ cw[53] ^ cw[55] ^ cw[57] ^ cw[59] ^ cw[61] ^ cw[63] ^ cw[65] ^ cw[67] ^ cw[69] ^ cw[71] ^ cw[73] ^ cw[74] ^ cw[77] ^ cw[79] ^ cw[81] ^ cw[83] ^ cw[85] ^ cw[86] ^ cw[89] ^ cw[91] ^ cw[93] ^ cw[95] ^ cw[97] ^ cw[98] ^ cw[100] ^ cw[102] ^ cw[104] ^ cw[106] ^ cw[109] ^ cw[111] ^ cw[113] ^ cw[115] ^ cw[117] ^ cw[119] ^ cw[121] ^ cw[123] ^ cw[125] ^ cw[127] ^ cw[128] ^ cw[131] ^ cw[133] ^ cw[135] ^ cw[137] ^ cw[139] ^ cw[140] ^ cw[142] ^ cw[144] ^ cw[146] ^ cw[148] ^ cw[151] ^ cw[153] ^ cw[155] ^ cw[157] ^ cw[159] ^ cw[161] ^ cw[163] ^ cw[165] ^ cw[167] ^ cw[169] ^ cw[170] ^ cw[172] ^ cw[174] ^ cw[176] ^ cw[178] ^ cw[181] ^ cw[183] ^ cw[185] ^ cw[187] ^ cw[189] ^ cw[191] ^ cw[193] ^ cw[195] ^ cw[197] ^ cw[199] ^ cw[200] ^ cw[202] ^ cw[204] ^ cw[206] ^ cw[208] ^ cw[210] ^ cw[212] ^ cw[214] ^ cw[216] ^ cw[218] ^ cw[221] ^ cw[223] ^ cw[225] ^ cw[227] ^ cw[229] ^ cw[231] ^ cw[233] ^ cw[235] ^ cw[237] ^ cw[239] ^ cw[240] ^ cw[243] ^ cw[245] ^ cw[247] ^ cw[249] ^ cw[251] ^ cw[252] ^ cw[254] ^ cw[256] ^ cw[258] ^ cw[260] ^ cw[263] ^ cw[265] ^ cw[267] ^ cw[269] ^ cw[271] ^ cw[273] ^ cw[275] ^ cw[277] ^ cw[279] ^ cw[281] ^ cw[282] ^ cw[284] ^ cw[286] ^ cw[288] ^ cw[290] ^ cw[293] ^ cw[295] ^ cw[297] ^ cw[299] ^ cw[301] ^ cw[303] ^ cw[305] ^ cw[307] ^ cw[309] ^ cw[311] ^ cw[312] ^ cw[314] ^ cw[316] ^ cw[318] ^ cw[320] ^ cw[322] ^ cw[324] ^ cw[326] ^ cw[328] ^ cw[330] ^ cw[333] ^ cw[335] ^ cw[337] ^ cw[339] ^ cw[341] ^ cw[343] ^ cw[345] ^ cw[347] ^ cw[349] ^ cw[351] ^ cw[352] ^ cw[354] ^ cw[356] ^ cw[358] ^ cw[360] ^ cw[363] ^ cw[365] ^ cw[367] ^ cw[369] ^ cw[371] ^ cw[373] ^ cw[375] ^ cw[377] ^ cw[379] ^ cw[381] ^ cw[382] ^ cw[384] ^ cw[386] ^ cw[388] ^ cw[390] ^ cw[392] ^ cw[394] ^ cw[396] ^ cw[398] ^ cw[400] ^ cw[403] ^ cw[405] ^ cw[407] ^ cw[409] ^ cw[411] ^ cw[413] ^ cw[415] ^ cw[417] ^ cw[419] ^ cw[421] ^ cw[422] ^ cw[424] ^ cw[426] ^ cw[428] ^ cw[430] ^ cw[432] ^ cw[434] ^ cw[436] ^ cw[438] ^ cw[440] ^ cw[443] ^ cw[445] ^ cw[447] ^ cw[449] ^ cw[451] ^ cw[453] ^ cw[455] ^ cw[457] ^ cw[459] ^ cw[461] ^ cw[462] ^ cw[464] ^ cw[466] ^ cw[468] ^ cw[470] ^ cw[472] ^ cw[474] ^ cw[476] ^ cw[478] ^ cw[480] ^ cw[483] ^ cw[485] ^ cw[487] ^ cw[489] ^ cw[491] ^ cw[492] ^ cw[493] ^ cw[494] ^ cw[495] ^ cw[496] ^ cw[498] ^ cw[499] ^ cw[500] ^ cw[501] ^ cw[507];
    assign syndrome[3] = cw[1] ^ cw[2] ^ cw[5] ^ cw[7] ^ cw[9] ^ cw[11] ^ cw[13] ^ cw[15] ^ cw[16] ^ cw[19] ^ cw[21] ^ cw[23] ^ cw[25] ^ cw[27] ^ cw[29] ^ cw[30] ^ cw[32] ^ cw[34] ^ cw[36] ^ cw[38] ^ cw[40] ^ cw[43] ^ cw[45] ^ cw[47] ^ cw[49] ^ cw[51] ^ cw[53] ^ cw[55] ^ cw[57] ^ cw[59] ^ cw[61] ^ cw[63] ^ cw[65] ^ cw[67] ^ cw[69] ^ cw[71] ^ cw[72] ^ cw[75] ^ cw[77] ^ cw[79] ^ cw[81] ^ cw[83] ^ cw[85] ^ cw[86] ^ cw[88] ^ cw[90] ^ cw[92] ^ cw[94] ^ cw[96] ^ cw[99] ^ cw[101] ^ cw[103] ^ cw[105] ^ cw[107] ^ cw[109] ^ cw[111] ^ cw[113] ^ cw[115] ^ cw[117] ^ cw[119] ^ cw[121] ^ cw[123] ^ cw[125] ^ cw[127] ^ cw[128] ^ cw[130] ^ cw[132] ^ cw[134] ^ cw[136] ^ cw[138] ^ cw[141] ^ cw[143] ^ cw[145] ^ cw[147] ^ cw[149] ^ cw[151] ^ cw[153] ^ cw[155] ^ cw[157] ^ cw[159] ^ cw[161] ^ cw[163] ^ cw[165] ^ cw[167] ^ cw[169] ^ cw[170] ^ cw[172] ^ cw[174] ^ cw[176] ^ cw[178] ^ cw[180] ^ cw[182] ^ cw[184] ^ cw[186] ^ cw[188] ^ cw[190] ^ cw[192] ^ cw[194] ^ cw[196] ^ cw[198] ^ cw[201] ^ cw[203] ^ cw[205] ^ cw[207] ^ cw[209] ^ cw[211] ^ cw[213] ^ cw[215] ^ cw[217] ^ cw[219] ^ cw[221] ^ cw[223] ^ cw[225] ^ cw[227] ^ cw[229] ^ cw[231] ^ cw[233] ^ cw[235] ^ cw[237] ^ cw[239] ^ cw[240] ^ cw[242] ^ cw[244] ^ cw[246] ^ cw[248] ^ cw[250] ^ cw[253] ^ cw[255] ^ cw[257] ^ cw[259] ^ cw[261] ^ cw[263] ^ cw[265] ^ cw[267] ^ cw[269] ^ cw[271] ^ cw[273] ^ cw[275] ^ cw[277] ^ cw[279] ^ cw[281] ^ cw[282] ^ cw[284] ^ cw[286] ^ cw[288] ^ cw[290] ^ cw[292] ^ cw[294] ^ cw[296] ^ cw[298] ^ cw[300] ^ cw[302] ^ cw[304] ^ cw[306] ^ cw[308] ^ cw[310] ^ cw[313] ^ cw[315] ^ cw[317] ^ cw[319] ^ cw[321] ^ cw[323] ^ cw[325] ^ cw[327] ^ cw[329] ^ cw[331] ^ cw[333] ^ cw[335] ^ cw[337] ^ cw[339] ^ cw[341] ^ cw[343] ^ cw[345] ^ cw[347] ^ cw[349] ^ cw[351] ^ cw[352] ^ cw[354] ^ cw[356] ^ cw[358] ^ cw[360] ^ cw[362] ^ cw[364] ^ cw[366] ^ cw[368] ^ cw[370] ^ cw[372] ^ cw[374] ^ cw[376] ^ cw[378] ^ cw[380] ^ cw[383] ^ cw[385] ^ cw[387] ^ cw[389] ^ cw[391] ^ cw[393] ^ cw[395] ^ cw[397] ^ cw[399] ^ cw[401] ^ cw[403] ^ cw[405] ^ cw[407] ^ cw[409] ^ cw[411] ^ cw[413] ^ cw[415] ^ cw[417] ^ cw[419] ^ cw[421] ^ cw[422] ^ cw[424] ^ cw[426] ^ cw[428] ^ cw[430] ^ cw[432] ^ cw[434] ^ cw[436] ^ cw[438] ^ cw[440] ^ cw[442] ^ cw[444] ^ cw[446] ^ cw[448] ^ cw[450] ^ cw[452] ^ cw[454] ^ cw[456] ^ cw[458] ^ cw[460] ^ cw[463] ^ cw[465] ^ cw[467] ^ cw[469] ^ cw[471] ^ cw[473] ^ cw[475] ^ cw[477] ^ cw[479] ^ cw[481] ^ cw[483] ^ cw[485] ^ cw[487] ^ cw[489] ^ cw[491] ^ cw[492] ^ cw[493] ^ cw[494] ^ cw[495] ^ cw[496] ^ cw[497] ^ cw[499] ^ cw[500] ^ cw[501] ^ cw[508];
    assign syndrome[2] = cw[0] ^ cw[3] ^ cw[5] ^ cw[7] ^ cw[9] ^ cw[11] ^ cw[13] ^ cw[15] ^ cw[16] ^ cw[18] ^ cw[20] ^ cw[22] ^ cw[24] ^ cw[26] ^ cw[28] ^ cw[31] ^ cw[33] ^ cw[35] ^ cw[37] ^ cw[39] ^ cw[41] ^ cw[43] ^ cw[45] ^ cw[47] ^ cw[49] ^ cw[51] ^ cw[53] ^ cw[55] ^ cw[57] ^ cw[59] ^ cw[61] ^ cw[63] ^ cw[65] ^ cw[67] ^ cw[69] ^ cw[71] ^ cw[72] ^ cw[74] ^ cw[76] ^ cw[78] ^ cw[80] ^ cw[82] ^ cw[84] ^ cw[87] ^ cw[89] ^ cw[91] ^ cw[93] ^ cw[95] ^ cw[97] ^ cw[99] ^ cw[101] ^ cw[103] ^ cw[105] ^ cw[107] ^ cw[109] ^ cw[111] ^ cw[113] ^ cw[115] ^ cw[117] ^ cw[119] ^ cw[121] ^ cw[123] ^ cw[125] ^ cw[127] ^ cw[128] ^ cw[130] ^ cw[132] ^ cw[134] ^ cw[136] ^ cw[138] ^ cw[140] ^ cw[142] ^ cw[144] ^ cw[146] ^ cw[148] ^ cw[150] ^ cw[152] ^ cw[154] ^ cw[156] ^ cw[158] ^ cw[160] ^ cw[162] ^ cw[164] ^ cw[166] ^ cw[168] ^ cw[171] ^ cw[173] ^ cw[175] ^ cw[177] ^ cw[179] ^ cw[181] ^ cw[183] ^ cw[185] ^ cw[187] ^ cw[189] ^ cw[191] ^ cw[193] ^ cw[195] ^ cw[197] ^ cw[199] ^ cw[201] ^ cw[203] ^ cw[205] ^ cw[207] ^ cw[209] ^ cw[211] ^ cw[213] ^ cw[215] ^ cw[217] ^ cw[219] ^ cw[221] ^ cw[223] ^ cw[225] ^ cw[227] ^ cw[229] ^ cw[231] ^ cw[233] ^ cw[235] ^ cw[237] ^ cw[239] ^ cw[240] ^ cw[242] ^ cw[244] ^ cw[246] ^ cw[248] ^ cw[250] ^ cw[252] ^ cw[254] ^ cw[256] ^ cw[258] ^ cw[260] ^ cw[262] ^ cw[264] ^ cw[266] ^ cw[268] ^ cw[270] ^ cw[272] ^ cw[274] ^ cw[276] ^ cw[278] ^ cw[280] ^ cw[283] ^ cw[285] ^ cw[287] ^ cw[289] ^ cw[291] ^ cw[293] ^ cw[295] ^ cw[297] ^ cw[299] ^ cw[301] ^ cw[303] ^ cw[305] ^ cw[307] ^ cw[309] ^ cw[311] ^ cw[313] ^ cw[315] ^ cw[317] ^ cw[319] ^ cw[321] ^ cw[323] ^ cw[325] ^ cw[327] ^ cw[329] ^ cw[331] ^ cw[333] ^ cw[335] ^ cw[337] ^ cw[339] ^ cw[341] ^ cw[343] ^ cw[345] ^ cw[347] ^ cw[349] ^ cw[351] ^ cw[352] ^ cw[354] ^ cw[356] ^ cw[358] ^ cw[360] ^ cw[362] ^ cw[364] ^ cw[366] ^ cw[368] ^ cw[370] ^ cw[372] ^ cw[374] ^ cw[376] ^ cw[378] ^ cw[380] ^ cw[382] ^ cw[384] ^ cw[386] ^ cw[388] ^ cw[390] ^ cw[392] ^ cw[394] ^ cw[396] ^ cw[398] ^ cw[400] ^ cw[402] ^ cw[404] ^ cw[406] ^ cw[408] ^ cw[410] ^ cw[412] ^ cw[414] ^ cw[416] ^ cw[418] ^ cw[420] ^ cw[423] ^ cw[425] ^ cw[427] ^ cw[429] ^ cw[431] ^ cw[433] ^ cw[435] ^ cw[437] ^ cw[439] ^ cw[441] ^ cw[443] ^ cw[445] ^ cw[447] ^ cw[449] ^ cw[451] ^ cw[453] ^ cw[455] ^ cw[457] ^ cw[459] ^ cw[461] ^ cw[463] ^ cw[465] ^ cw[467] ^ cw[469] ^ cw[471] ^ cw[473] ^ cw[475] ^ cw[477] ^ cw[479] ^ cw[481] ^ cw[483] ^ cw[485] ^ cw[487] ^ cw[489] ^ cw[491] ^ cw[492] ^ cw[493] ^ cw[494] ^ cw[495] ^ cw[496] ^ cw[497] ^ cw[498] ^ cw[500] ^ cw[501] ^ cw[509];
    assign syndrome[1] = cw[0] ^ cw[2] ^ cw[4] ^ cw[6] ^ cw[8] ^ cw[10] ^ cw[12] ^ cw[14] ^ cw[17] ^ cw[19] ^ cw[21] ^ cw[23] ^ cw[25] ^ cw[27] ^ cw[29] ^ cw[31] ^ cw[33] ^ cw[35] ^ cw[37] ^ cw[39] ^ cw[41] ^ cw[43] ^ cw[45] ^ cw[47] ^ cw[49] ^ cw[51] ^ cw[53] ^ cw[55] ^ cw[57] ^ cw[59] ^ cw[61] ^ cw[63] ^ cw[65] ^ cw[67] ^ cw[69] ^ cw[71] ^ cw[72] ^ cw[74] ^ cw[76] ^ cw[78] ^ cw[80] ^ cw[82] ^ cw[84] ^ cw[86] ^ cw[88] ^ cw[90] ^ cw[92] ^ cw[94] ^ cw[96] ^ cw[98] ^ cw[100] ^ cw[102] ^ cw[104] ^ cw[106] ^ cw[108] ^ cw[110] ^ cw[112] ^ cw[114] ^ cw[116] ^ cw[118] ^ cw[120] ^ cw[122] ^ cw[124] ^ cw[126] ^ cw[129] ^ cw[131] ^ cw[133] ^ cw[135] ^ cw[137] ^ cw[139] ^ cw[141] ^ cw[143] ^ cw[145] ^ cw[147] ^ cw[149] ^ cw[151] ^ cw[153] ^ cw[155] ^ cw[157] ^ cw[159] ^ cw[161] ^ cw[163] ^ cw[165] ^ cw[167] ^ cw[169] ^ cw[171] ^ cw[173] ^ cw[175] ^ cw[177] ^ cw[179] ^ cw[181] ^ cw[183] ^ cw[185] ^ cw[187] ^ cw[189] ^ cw[191] ^ cw[193] ^ cw[195] ^ cw[197] ^ cw[199] ^ cw[201] ^ cw[203] ^ cw[205] ^ cw[207] ^ cw[209] ^ cw[211] ^ cw[213] ^ cw[215] ^ cw[217] ^ cw[219] ^ cw[221] ^ cw[223] ^ cw[225] ^ cw[227] ^ cw[229] ^ cw[231] ^ cw[233] ^ cw[235] ^ cw[237] ^ cw[239] ^ cw[240] ^ cw[242] ^ cw[244] ^ cw[246] ^ cw[248] ^ cw[250] ^ cw[252] ^ cw[254] ^ cw[256] ^ cw[258] ^ cw[260] ^ cw[262] ^ cw[264] ^ cw[266] ^ cw[268] ^ cw[270] ^ cw[272] ^ cw[274] ^ cw[276] ^ cw[278] ^ cw[280] ^ cw[282] ^ cw[284] ^ cw[286] ^ cw[288] ^ cw[290] ^ cw[292] ^ cw[294] ^ cw[296] ^ cw[298] ^ cw[300] ^ cw[302] ^ cw[304] ^ cw[306] ^ cw[308] ^ cw[310] ^ cw[312] ^ cw[314] ^ cw[316] ^ cw[318] ^ cw[320] ^ cw[322] ^ cw[324] ^ cw[326] ^ cw[328] ^ cw[330] ^ cw[332] ^ cw[334] ^ cw[336] ^ cw[338] ^ cw[340] ^ cw[342] ^ cw[344] ^ cw[346] ^ cw[348] ^ cw[350] ^ cw[353] ^ cw[355] ^ cw[357] ^ cw[359] ^ cw[361] ^ cw[363] ^ cw[365] ^ cw[367] ^ cw[369] ^ cw[371] ^ cw[373] ^ cw[375] ^ cw[377] ^ cw[379] ^ cw[381] ^ cw[383] ^ cw[385] ^ cw[387] ^ cw[389] ^ cw[391] ^ cw[393] ^ cw[395] ^ cw[397] ^ cw[399] ^ cw[401] ^ cw[403] ^ cw[405] ^ cw[407] ^ cw[409] ^ cw[411] ^ cw[413] ^ cw[415] ^ cw[417] ^ cw[419] ^ cw[421] ^ cw[423] ^ cw[425] ^ cw[427] ^ cw[429] ^ cw[431] ^ cw[433] ^ cw[435] ^ cw[437] ^ cw[439] ^ cw[441] ^ cw[443] ^ cw[445] ^ cw[447] ^ cw[449] ^ cw[451] ^ cw[453] ^ cw[455] ^ cw[457] ^ cw[459] ^ cw[461] ^ cw[463] ^ cw[465] ^ cw[467] ^ cw[469] ^ cw[471] ^ cw[473] ^ cw[475] ^ cw[477] ^ cw[479] ^ cw[481] ^ cw[483] ^ cw[485] ^ cw[487] ^ cw[489] ^ cw[491] ^ cw[492] ^ cw[493] ^ cw[494] ^ cw[495] ^ cw[496] ^ cw[497] ^ cw[498] ^ cw[499] ^ cw[501] ^ cw[510];
    assign syndrome[0] = cw[0] ^ cw[2] ^ cw[4] ^ cw[6] ^ cw[8] ^ cw[10] ^ cw[12] ^ cw[14] ^ cw[16] ^ cw[18] ^ cw[20] ^ cw[22] ^ cw[24] ^ cw[26] ^ cw[28] ^ cw[30] ^ cw[32] ^ cw[34] ^ cw[36] ^ cw[38] ^ cw[40] ^ cw[42] ^ cw[44] ^ cw[46] ^ cw[48] ^ cw[50] ^ cw[52] ^ cw[54] ^ cw[56] ^ cw[58] ^ cw[60] ^ cw[62] ^ cw[64] ^ cw[66] ^ cw[68] ^ cw[70] ^ cw[73] ^ cw[75] ^ cw[77] ^ cw[79] ^ cw[81] ^ cw[83] ^ cw[85] ^ cw[87] ^ cw[89] ^ cw[91] ^ cw[93] ^ cw[95] ^ cw[97] ^ cw[99] ^ cw[101] ^ cw[103] ^ cw[105] ^ cw[107] ^ cw[109] ^ cw[111] ^ cw[113] ^ cw[115] ^ cw[117] ^ cw[119] ^ cw[121] ^ cw[123] ^ cw[125] ^ cw[127] ^ cw[129] ^ cw[131] ^ cw[133] ^ cw[135] ^ cw[137] ^ cw[139] ^ cw[141] ^ cw[143] ^ cw[145] ^ cw[147] ^ cw[149] ^ cw[151] ^ cw[153] ^ cw[155] ^ cw[157] ^ cw[159] ^ cw[161] ^ cw[163] ^ cw[165] ^ cw[167] ^ cw[169] ^ cw[171] ^ cw[173] ^ cw[175] ^ cw[177] ^ cw[179] ^ cw[181] ^ cw[183] ^ cw[185] ^ cw[187] ^ cw[189] ^ cw[191] ^ cw[193] ^ cw[195] ^ cw[197] ^ cw[199] ^ cw[201] ^ cw[203] ^ cw[205] ^ cw[207] ^ cw[209] ^ cw[211] ^ cw[213] ^ cw[215] ^ cw[217] ^ cw[219] ^ cw[221] ^ cw[223] ^ cw[225] ^ cw[227] ^ cw[229] ^ cw[231] ^ cw[233] ^ cw[235] ^ cw[237] ^ cw[239] ^ cw[240] ^ cw[242] ^ cw[244] ^ cw[246] ^ cw[248] ^ cw[250] ^ cw[252] ^ cw[254] ^ cw[256] ^ cw[258] ^ cw[260] ^ cw[262] ^ cw[264] ^ cw[266] ^ cw[268] ^ cw[270] ^ cw[272] ^ cw[274] ^ cw[276] ^ cw[278] ^ cw[280] ^ cw[282] ^ cw[284] ^ cw[286] ^ cw[288] ^ cw[290] ^ cw[292] ^ cw[294] ^ cw[296] ^ cw[298] ^ cw[300] ^ cw[302] ^ cw[304] ^ cw[306] ^ cw[308] ^ cw[310] ^ cw[312] ^ cw[314] ^ cw[316] ^ cw[318] ^ cw[320] ^ cw[322] ^ cw[324] ^ cw[326] ^ cw[328] ^ cw[330] ^ cw[332] ^ cw[334] ^ cw[336] ^ cw[338] ^ cw[340] ^ cw[342] ^ cw[344] ^ cw[346] ^ cw[348] ^ cw[350] ^ cw[352] ^ cw[354] ^ cw[356] ^ cw[358] ^ cw[360] ^ cw[362] ^ cw[364] ^ cw[366] ^ cw[368] ^ cw[370] ^ cw[372] ^ cw[374] ^ cw[376] ^ cw[378] ^ cw[380] ^ cw[382] ^ cw[384] ^ cw[386] ^ cw[388] ^ cw[390] ^ cw[392] ^ cw[394] ^ cw[396] ^ cw[398] ^ cw[400] ^ cw[402] ^ cw[404] ^ cw[406] ^ cw[408] ^ cw[410] ^ cw[412] ^ cw[414] ^ cw[416] ^ cw[418] ^ cw[420] ^ cw[422] ^ cw[424] ^ cw[426] ^ cw[428] ^ cw[430] ^ cw[432] ^ cw[434] ^ cw[436] ^ cw[438] ^ cw[440] ^ cw[442] ^ cw[444] ^ cw[446] ^ cw[448] ^ cw[450] ^ cw[452] ^ cw[454] ^ cw[456] ^ cw[458] ^ cw[460] ^ cw[462] ^ cw[464] ^ cw[466] ^ cw[468] ^ cw[470] ^ cw[472] ^ cw[474] ^ cw[476] ^ cw[478] ^ cw[480] ^ cw[482] ^ cw[484] ^ cw[486] ^ cw[488] ^ cw[490] ^ cw[492] ^ cw[493] ^ cw[494] ^ cw[495] ^ cw[496] ^ cw[497] ^ cw[498] ^ cw[499] ^ cw[500] ^ cw[511];
    assign parity_check_matrix[0] = 10'b0000000111;
    assign parity_check_matrix[1] = 10'b1111111000;
    assign parity_check_matrix[2] = 10'b0000001011;
    assign parity_check_matrix[3] = 10'b1111110100;
    assign parity_check_matrix[4] = 10'b0000010011;
    assign parity_check_matrix[5] = 10'b1111101100;
    assign parity_check_matrix[6] = 10'b0000100011;
    assign parity_check_matrix[7] = 10'b1111011100;
    assign parity_check_matrix[8] = 10'b0001000011;
    assign parity_check_matrix[9] = 10'b1110111100;
    assign parity_check_matrix[10] = 10'b0010000011;
    assign parity_check_matrix[11] = 10'b1101111100;
    assign parity_check_matrix[12] = 10'b0100000011;
    assign parity_check_matrix[13] = 10'b1011111100;
    assign parity_check_matrix[14] = 10'b1000000011;
    assign parity_check_matrix[15] = 10'b0111111100;
    assign parity_check_matrix[16] = 10'b0000001101;
    assign parity_check_matrix[17] = 10'b1111110010;
    assign parity_check_matrix[18] = 10'b0000010101;
    assign parity_check_matrix[19] = 10'b1111101010;
    assign parity_check_matrix[20] = 10'b0000100101;
    assign parity_check_matrix[21] = 10'b1111011010;
    assign parity_check_matrix[22] = 10'b0001000101;
    assign parity_check_matrix[23] = 10'b1110111010;
    assign parity_check_matrix[24] = 10'b0010000101;
    assign parity_check_matrix[25] = 10'b1101111010;
    assign parity_check_matrix[26] = 10'b0100000101;
    assign parity_check_matrix[27] = 10'b1011111010;
    assign parity_check_matrix[28] = 10'b1000000101;
    assign parity_check_matrix[29] = 10'b0111111010;
    assign parity_check_matrix[30] = 10'b0000011001;
    assign parity_check_matrix[31] = 10'b1111100110;
    assign parity_check_matrix[32] = 10'b0000101001;
    assign parity_check_matrix[33] = 10'b1111010110;
    assign parity_check_matrix[34] = 10'b0001001001;
    assign parity_check_matrix[35] = 10'b1110110110;
    assign parity_check_matrix[36] = 10'b0010001001;
    assign parity_check_matrix[37] = 10'b1101110110;
    assign parity_check_matrix[38] = 10'b0100001001;
    assign parity_check_matrix[39] = 10'b1011110110;
    assign parity_check_matrix[40] = 10'b1000001001;
    assign parity_check_matrix[41] = 10'b0111110110;
    assign parity_check_matrix[42] = 10'b0000110001;
    assign parity_check_matrix[43] = 10'b1111001110;
    assign parity_check_matrix[44] = 10'b0001010001;
    assign parity_check_matrix[45] = 10'b1110101110;
    assign parity_check_matrix[46] = 10'b0010010001;
    assign parity_check_matrix[47] = 10'b1101101110;
    assign parity_check_matrix[48] = 10'b0100010001;
    assign parity_check_matrix[49] = 10'b1011101110;
    assign parity_check_matrix[50] = 10'b1000010001;
    assign parity_check_matrix[51] = 10'b0111101110;
    assign parity_check_matrix[52] = 10'b0001100001;
    assign parity_check_matrix[53] = 10'b1110011110;
    assign parity_check_matrix[54] = 10'b0010100001;
    assign parity_check_matrix[55] = 10'b1101011110;
    assign parity_check_matrix[56] = 10'b0100100001;
    assign parity_check_matrix[57] = 10'b1011011110;
    assign parity_check_matrix[58] = 10'b1000100001;
    assign parity_check_matrix[59] = 10'b0111011110;
    assign parity_check_matrix[60] = 10'b0011000001;
    assign parity_check_matrix[61] = 10'b1100111110;
    assign parity_check_matrix[62] = 10'b0101000001;
    assign parity_check_matrix[63] = 10'b1010111110;
    assign parity_check_matrix[64] = 10'b1001000001;
    assign parity_check_matrix[65] = 10'b0110111110;
    assign parity_check_matrix[66] = 10'b0110000001;
    assign parity_check_matrix[67] = 10'b1001111110;
    assign parity_check_matrix[68] = 10'b1010000001;
    assign parity_check_matrix[69] = 10'b0101111110;
    assign parity_check_matrix[70] = 10'b1100000001;
    assign parity_check_matrix[71] = 10'b0011111110;
    assign parity_check_matrix[72] = 10'b0000001110;
    assign parity_check_matrix[73] = 10'b1111110001;
    assign parity_check_matrix[74] = 10'b0000010110;
    assign parity_check_matrix[75] = 10'b1111101001;
    assign parity_check_matrix[76] = 10'b0000100110;
    assign parity_check_matrix[77] = 10'b1111011001;
    assign parity_check_matrix[78] = 10'b0001000110;
    assign parity_check_matrix[79] = 10'b1110111001;
    assign parity_check_matrix[80] = 10'b0010000110;
    assign parity_check_matrix[81] = 10'b1101111001;
    assign parity_check_matrix[82] = 10'b0100000110;
    assign parity_check_matrix[83] = 10'b1011111001;
    assign parity_check_matrix[84] = 10'b1000000110;
    assign parity_check_matrix[85] = 10'b0111111001;
    assign parity_check_matrix[86] = 10'b0000011010;
    assign parity_check_matrix[87] = 10'b1111100101;
    assign parity_check_matrix[88] = 10'b0000101010;
    assign parity_check_matrix[89] = 10'b1111010101;
    assign parity_check_matrix[90] = 10'b0001001010;
    assign parity_check_matrix[91] = 10'b1110110101;
    assign parity_check_matrix[92] = 10'b0010001010;
    assign parity_check_matrix[93] = 10'b1101110101;
    assign parity_check_matrix[94] = 10'b0100001010;
    assign parity_check_matrix[95] = 10'b1011110101;
    assign parity_check_matrix[96] = 10'b1000001010;
    assign parity_check_matrix[97] = 10'b0111110101;
    assign parity_check_matrix[98] = 10'b0000110010;
    assign parity_check_matrix[99] = 10'b1111001101;
    assign parity_check_matrix[100] = 10'b0001010010;
    assign parity_check_matrix[101] = 10'b1110101101;
    assign parity_check_matrix[102] = 10'b0010010010;
    assign parity_check_matrix[103] = 10'b1101101101;
    assign parity_check_matrix[104] = 10'b0100010010;
    assign parity_check_matrix[105] = 10'b1011101101;
    assign parity_check_matrix[106] = 10'b1000010010;
    assign parity_check_matrix[107] = 10'b0111101101;
    assign parity_check_matrix[108] = 10'b0001100010;
    assign parity_check_matrix[109] = 10'b1110011101;
    assign parity_check_matrix[110] = 10'b0010100010;
    assign parity_check_matrix[111] = 10'b1101011101;
    assign parity_check_matrix[112] = 10'b0100100010;
    assign parity_check_matrix[113] = 10'b1011011101;
    assign parity_check_matrix[114] = 10'b1000100010;
    assign parity_check_matrix[115] = 10'b0111011101;
    assign parity_check_matrix[116] = 10'b0011000010;
    assign parity_check_matrix[117] = 10'b1100111101;
    assign parity_check_matrix[118] = 10'b0101000010;
    assign parity_check_matrix[119] = 10'b1010111101;
    assign parity_check_matrix[120] = 10'b1001000010;
    assign parity_check_matrix[121] = 10'b0110111101;
    assign parity_check_matrix[122] = 10'b0110000010;
    assign parity_check_matrix[123] = 10'b1001111101;
    assign parity_check_matrix[124] = 10'b1010000010;
    assign parity_check_matrix[125] = 10'b0101111101;
    assign parity_check_matrix[126] = 10'b1100000010;
    assign parity_check_matrix[127] = 10'b0011111101;
    assign parity_check_matrix[128] = 10'b0000011100;
    assign parity_check_matrix[129] = 10'b1111100011;
    assign parity_check_matrix[130] = 10'b0000101100;
    assign parity_check_matrix[131] = 10'b1111010011;
    assign parity_check_matrix[132] = 10'b0001001100;
    assign parity_check_matrix[133] = 10'b1110110011;
    assign parity_check_matrix[134] = 10'b0010001100;
    assign parity_check_matrix[135] = 10'b1101110011;
    assign parity_check_matrix[136] = 10'b0100001100;
    assign parity_check_matrix[137] = 10'b1011110011;
    assign parity_check_matrix[138] = 10'b1000001100;
    assign parity_check_matrix[139] = 10'b0111110011;
    assign parity_check_matrix[140] = 10'b0000110100;
    assign parity_check_matrix[141] = 10'b1111001011;
    assign parity_check_matrix[142] = 10'b0001010100;
    assign parity_check_matrix[143] = 10'b1110101011;
    assign parity_check_matrix[144] = 10'b0010010100;
    assign parity_check_matrix[145] = 10'b1101101011;
    assign parity_check_matrix[146] = 10'b0100010100;
    assign parity_check_matrix[147] = 10'b1011101011;
    assign parity_check_matrix[148] = 10'b1000010100;
    assign parity_check_matrix[149] = 10'b0111101011;
    assign parity_check_matrix[150] = 10'b0001100100;
    assign parity_check_matrix[151] = 10'b1110011011;
    assign parity_check_matrix[152] = 10'b0010100100;
    assign parity_check_matrix[153] = 10'b1101011011;
    assign parity_check_matrix[154] = 10'b0100100100;
    assign parity_check_matrix[155] = 10'b1011011011;
    assign parity_check_matrix[156] = 10'b1000100100;
    assign parity_check_matrix[157] = 10'b0111011011;
    assign parity_check_matrix[158] = 10'b0011000100;
    assign parity_check_matrix[159] = 10'b1100111011;
    assign parity_check_matrix[160] = 10'b0101000100;
    assign parity_check_matrix[161] = 10'b1010111011;
    assign parity_check_matrix[162] = 10'b1001000100;
    assign parity_check_matrix[163] = 10'b0110111011;
    assign parity_check_matrix[164] = 10'b0110000100;
    assign parity_check_matrix[165] = 10'b1001111011;
    assign parity_check_matrix[166] = 10'b1010000100;
    assign parity_check_matrix[167] = 10'b0101111011;
    assign parity_check_matrix[168] = 10'b1100000100;
    assign parity_check_matrix[169] = 10'b0011111011;
    assign parity_check_matrix[170] = 10'b0000111000;
    assign parity_check_matrix[171] = 10'b1111000111;
    assign parity_check_matrix[172] = 10'b0001011000;
    assign parity_check_matrix[173] = 10'b1110100111;
    assign parity_check_matrix[174] = 10'b0010011000;
    assign parity_check_matrix[175] = 10'b1101100111;
    assign parity_check_matrix[176] = 10'b0100011000;
    assign parity_check_matrix[177] = 10'b1011100111;
    assign parity_check_matrix[178] = 10'b1000011000;
    assign parity_check_matrix[179] = 10'b0111100111;
    assign parity_check_matrix[180] = 10'b0001101000;
    assign parity_check_matrix[181] = 10'b1110010111;
    assign parity_check_matrix[182] = 10'b0010101000;
    assign parity_check_matrix[183] = 10'b1101010111;
    assign parity_check_matrix[184] = 10'b0100101000;
    assign parity_check_matrix[185] = 10'b1011010111;
    assign parity_check_matrix[186] = 10'b1000101000;
    assign parity_check_matrix[187] = 10'b0111010111;
    assign parity_check_matrix[188] = 10'b0011001000;
    assign parity_check_matrix[189] = 10'b1100110111;
    assign parity_check_matrix[190] = 10'b0101001000;
    assign parity_check_matrix[191] = 10'b1010110111;
    assign parity_check_matrix[192] = 10'b1001001000;
    assign parity_check_matrix[193] = 10'b0110110111;
    assign parity_check_matrix[194] = 10'b0110001000;
    assign parity_check_matrix[195] = 10'b1001110111;
    assign parity_check_matrix[196] = 10'b1010001000;
    assign parity_check_matrix[197] = 10'b0101110111;
    assign parity_check_matrix[198] = 10'b1100001000;
    assign parity_check_matrix[199] = 10'b0011110111;
    assign parity_check_matrix[200] = 10'b0001110000;
    assign parity_check_matrix[201] = 10'b1110001111;
    assign parity_check_matrix[202] = 10'b0010110000;
    assign parity_check_matrix[203] = 10'b1101001111;
    assign parity_check_matrix[204] = 10'b0100110000;
    assign parity_check_matrix[205] = 10'b1011001111;
    assign parity_check_matrix[206] = 10'b1000110000;
    assign parity_check_matrix[207] = 10'b0111001111;
    assign parity_check_matrix[208] = 10'b0011010000;
    assign parity_check_matrix[209] = 10'b1100101111;
    assign parity_check_matrix[210] = 10'b0101010000;
    assign parity_check_matrix[211] = 10'b1010101111;
    assign parity_check_matrix[212] = 10'b1001010000;
    assign parity_check_matrix[213] = 10'b0110101111;
    assign parity_check_matrix[214] = 10'b0110010000;
    assign parity_check_matrix[215] = 10'b1001101111;
    assign parity_check_matrix[216] = 10'b1010010000;
    assign parity_check_matrix[217] = 10'b0101101111;
    assign parity_check_matrix[218] = 10'b1100010000;
    assign parity_check_matrix[219] = 10'b0011101111;
    assign parity_check_matrix[220] = 10'b0011100000;
    assign parity_check_matrix[221] = 10'b1100011111;
    assign parity_check_matrix[222] = 10'b0101100000;
    assign parity_check_matrix[223] = 10'b1010011111;
    assign parity_check_matrix[224] = 10'b1001100000;
    assign parity_check_matrix[225] = 10'b0110011111;
    assign parity_check_matrix[226] = 10'b0110100000;
    assign parity_check_matrix[227] = 10'b1001011111;
    assign parity_check_matrix[228] = 10'b1010100000;
    assign parity_check_matrix[229] = 10'b0101011111;
    assign parity_check_matrix[230] = 10'b1100100000;
    assign parity_check_matrix[231] = 10'b0011011111;
    assign parity_check_matrix[232] = 10'b0111000000;
    assign parity_check_matrix[233] = 10'b1000111111;
    assign parity_check_matrix[234] = 10'b1011000000;
    assign parity_check_matrix[235] = 10'b0100111111;
    assign parity_check_matrix[236] = 10'b1101000000;
    assign parity_check_matrix[237] = 10'b0010111111;
    assign parity_check_matrix[238] = 10'b1110000000;
    assign parity_check_matrix[239] = 10'b0001111111;
    assign parity_check_matrix[240] = 10'b0000011111;
    assign parity_check_matrix[241] = 10'b1111100000;
    assign parity_check_matrix[242] = 10'b0000101111;
    assign parity_check_matrix[243] = 10'b1111010000;
    assign parity_check_matrix[244] = 10'b0001001111;
    assign parity_check_matrix[245] = 10'b1110110000;
    assign parity_check_matrix[246] = 10'b0010001111;
    assign parity_check_matrix[247] = 10'b1101110000;
    assign parity_check_matrix[248] = 10'b0100001111;
    assign parity_check_matrix[249] = 10'b1011110000;
    assign parity_check_matrix[250] = 10'b1000001111;
    assign parity_check_matrix[251] = 10'b0111110000;
    assign parity_check_matrix[252] = 10'b0000110111;
    assign parity_check_matrix[253] = 10'b1111001000;
    assign parity_check_matrix[254] = 10'b0001010111;
    assign parity_check_matrix[255] = 10'b1110101000;
    assign parity_check_matrix[256] = 10'b0010010111;
    assign parity_check_matrix[257] = 10'b1101101000;
    assign parity_check_matrix[258] = 10'b0100010111;
    assign parity_check_matrix[259] = 10'b1011101000;
    assign parity_check_matrix[260] = 10'b1000010111;
    assign parity_check_matrix[261] = 10'b0111101000;
    assign parity_check_matrix[262] = 10'b0001100111;
    assign parity_check_matrix[263] = 10'b1110011000;
    assign parity_check_matrix[264] = 10'b0010100111;
    assign parity_check_matrix[265] = 10'b1101011000;
    assign parity_check_matrix[266] = 10'b0100100111;
    assign parity_check_matrix[267] = 10'b1011011000;
    assign parity_check_matrix[268] = 10'b1000100111;
    assign parity_check_matrix[269] = 10'b0111011000;
    assign parity_check_matrix[270] = 10'b0011000111;
    assign parity_check_matrix[271] = 10'b1100111000;
    assign parity_check_matrix[272] = 10'b0101000111;
    assign parity_check_matrix[273] = 10'b1010111000;
    assign parity_check_matrix[274] = 10'b1001000111;
    assign parity_check_matrix[275] = 10'b0110111000;
    assign parity_check_matrix[276] = 10'b0110000111;
    assign parity_check_matrix[277] = 10'b1001111000;
    assign parity_check_matrix[278] = 10'b1010000111;
    assign parity_check_matrix[279] = 10'b0101111000;
    assign parity_check_matrix[280] = 10'b1100000111;
    assign parity_check_matrix[281] = 10'b0011111000;
    assign parity_check_matrix[282] = 10'b0000111011;
    assign parity_check_matrix[283] = 10'b1111000100;
    assign parity_check_matrix[284] = 10'b0001011011;
    assign parity_check_matrix[285] = 10'b1110100100;
    assign parity_check_matrix[286] = 10'b0010011011;
    assign parity_check_matrix[287] = 10'b1101100100;
    assign parity_check_matrix[288] = 10'b0100011011;
    assign parity_check_matrix[289] = 10'b1011100100;
    assign parity_check_matrix[290] = 10'b1000011011;
    assign parity_check_matrix[291] = 10'b0111100100;
    assign parity_check_matrix[292] = 10'b0001101011;
    assign parity_check_matrix[293] = 10'b1110010100;
    assign parity_check_matrix[294] = 10'b0010101011;
    assign parity_check_matrix[295] = 10'b1101010100;
    assign parity_check_matrix[296] = 10'b0100101011;
    assign parity_check_matrix[297] = 10'b1011010100;
    assign parity_check_matrix[298] = 10'b1000101011;
    assign parity_check_matrix[299] = 10'b0111010100;
    assign parity_check_matrix[300] = 10'b0011001011;
    assign parity_check_matrix[301] = 10'b1100110100;
    assign parity_check_matrix[302] = 10'b0101001011;
    assign parity_check_matrix[303] = 10'b1010110100;
    assign parity_check_matrix[304] = 10'b1001001011;
    assign parity_check_matrix[305] = 10'b0110110100;
    assign parity_check_matrix[306] = 10'b0110001011;
    assign parity_check_matrix[307] = 10'b1001110100;
    assign parity_check_matrix[308] = 10'b1010001011;
    assign parity_check_matrix[309] = 10'b0101110100;
    assign parity_check_matrix[310] = 10'b1100001011;
    assign parity_check_matrix[311] = 10'b0011110100;
    assign parity_check_matrix[312] = 10'b0001110011;
    assign parity_check_matrix[313] = 10'b1110001100;
    assign parity_check_matrix[314] = 10'b0010110011;
    assign parity_check_matrix[315] = 10'b1101001100;
    assign parity_check_matrix[316] = 10'b0100110011;
    assign parity_check_matrix[317] = 10'b1011001100;
    assign parity_check_matrix[318] = 10'b1000110011;
    assign parity_check_matrix[319] = 10'b0111001100;
    assign parity_check_matrix[320] = 10'b0011010011;
    assign parity_check_matrix[321] = 10'b1100101100;
    assign parity_check_matrix[322] = 10'b0101010011;
    assign parity_check_matrix[323] = 10'b1010101100;
    assign parity_check_matrix[324] = 10'b1001010011;
    assign parity_check_matrix[325] = 10'b0110101100;
    assign parity_check_matrix[326] = 10'b0110010011;
    assign parity_check_matrix[327] = 10'b1001101100;
    assign parity_check_matrix[328] = 10'b1010010011;
    assign parity_check_matrix[329] = 10'b0101101100;
    assign parity_check_matrix[330] = 10'b1100010011;
    assign parity_check_matrix[331] = 10'b0011101100;
    assign parity_check_matrix[332] = 10'b0011100011;
    assign parity_check_matrix[333] = 10'b1100011100;
    assign parity_check_matrix[334] = 10'b0101100011;
    assign parity_check_matrix[335] = 10'b1010011100;
    assign parity_check_matrix[336] = 10'b1001100011;
    assign parity_check_matrix[337] = 10'b0110011100;
    assign parity_check_matrix[338] = 10'b0110100011;
    assign parity_check_matrix[339] = 10'b1001011100;
    assign parity_check_matrix[340] = 10'b1010100011;
    assign parity_check_matrix[341] = 10'b0101011100;
    assign parity_check_matrix[342] = 10'b1100100011;
    assign parity_check_matrix[343] = 10'b0011011100;
    assign parity_check_matrix[344] = 10'b0111000011;
    assign parity_check_matrix[345] = 10'b1000111100;
    assign parity_check_matrix[346] = 10'b1011000011;
    assign parity_check_matrix[347] = 10'b0100111100;
    assign parity_check_matrix[348] = 10'b1101000011;
    assign parity_check_matrix[349] = 10'b0010111100;
    assign parity_check_matrix[350] = 10'b1110000011;
    assign parity_check_matrix[351] = 10'b0001111100;
    assign parity_check_matrix[352] = 10'b0000111101;
    assign parity_check_matrix[353] = 10'b1111000010;
    assign parity_check_matrix[354] = 10'b0001011101;
    assign parity_check_matrix[355] = 10'b1110100010;
    assign parity_check_matrix[356] = 10'b0010011101;
    assign parity_check_matrix[357] = 10'b1101100010;
    assign parity_check_matrix[358] = 10'b0100011101;
    assign parity_check_matrix[359] = 10'b1011100010;
    assign parity_check_matrix[360] = 10'b1000011101;
    assign parity_check_matrix[361] = 10'b0111100010;
    assign parity_check_matrix[362] = 10'b0001101101;
    assign parity_check_matrix[363] = 10'b1110010010;
    assign parity_check_matrix[364] = 10'b0010101101;
    assign parity_check_matrix[365] = 10'b1101010010;
    assign parity_check_matrix[366] = 10'b0100101101;
    assign parity_check_matrix[367] = 10'b1011010010;
    assign parity_check_matrix[368] = 10'b1000101101;
    assign parity_check_matrix[369] = 10'b0111010010;
    assign parity_check_matrix[370] = 10'b0011001101;
    assign parity_check_matrix[371] = 10'b1100110010;
    assign parity_check_matrix[372] = 10'b0101001101;
    assign parity_check_matrix[373] = 10'b1010110010;
    assign parity_check_matrix[374] = 10'b1001001101;
    assign parity_check_matrix[375] = 10'b0110110010;
    assign parity_check_matrix[376] = 10'b0110001101;
    assign parity_check_matrix[377] = 10'b1001110010;
    assign parity_check_matrix[378] = 10'b1010001101;
    assign parity_check_matrix[379] = 10'b0101110010;
    assign parity_check_matrix[380] = 10'b1100001101;
    assign parity_check_matrix[381] = 10'b0011110010;
    assign parity_check_matrix[382] = 10'b0001110101;
    assign parity_check_matrix[383] = 10'b1110001010;
    assign parity_check_matrix[384] = 10'b0010110101;
    assign parity_check_matrix[385] = 10'b1101001010;
    assign parity_check_matrix[386] = 10'b0100110101;
    assign parity_check_matrix[387] = 10'b1011001010;
    assign parity_check_matrix[388] = 10'b1000110101;
    assign parity_check_matrix[389] = 10'b0111001010;
    assign parity_check_matrix[390] = 10'b0011010101;
    assign parity_check_matrix[391] = 10'b1100101010;
    assign parity_check_matrix[392] = 10'b0101010101;
    assign parity_check_matrix[393] = 10'b1010101010;
    assign parity_check_matrix[394] = 10'b1001010101;
    assign parity_check_matrix[395] = 10'b0110101010;
    assign parity_check_matrix[396] = 10'b0110010101;
    assign parity_check_matrix[397] = 10'b1001101010;
    assign parity_check_matrix[398] = 10'b1010010101;
    assign parity_check_matrix[399] = 10'b0101101010;
    assign parity_check_matrix[400] = 10'b1100010101;
    assign parity_check_matrix[401] = 10'b0011101010;
    assign parity_check_matrix[402] = 10'b0011100101;
    assign parity_check_matrix[403] = 10'b1100011010;
    assign parity_check_matrix[404] = 10'b0101100101;
    assign parity_check_matrix[405] = 10'b1010011010;
    assign parity_check_matrix[406] = 10'b1001100101;
    assign parity_check_matrix[407] = 10'b0110011010;
    assign parity_check_matrix[408] = 10'b0110100101;
    assign parity_check_matrix[409] = 10'b1001011010;
    assign parity_check_matrix[410] = 10'b1010100101;
    assign parity_check_matrix[411] = 10'b0101011010;
    assign parity_check_matrix[412] = 10'b1100100101;
    assign parity_check_matrix[413] = 10'b0011011010;
    assign parity_check_matrix[414] = 10'b0111000101;
    assign parity_check_matrix[415] = 10'b1000111010;
    assign parity_check_matrix[416] = 10'b1011000101;
    assign parity_check_matrix[417] = 10'b0100111010;
    assign parity_check_matrix[418] = 10'b1101000101;
    assign parity_check_matrix[419] = 10'b0010111010;
    assign parity_check_matrix[420] = 10'b1110000101;
    assign parity_check_matrix[421] = 10'b0001111010;
    assign parity_check_matrix[422] = 10'b0001111001;
    assign parity_check_matrix[423] = 10'b1110000110;
    assign parity_check_matrix[424] = 10'b0010111001;
    assign parity_check_matrix[425] = 10'b1101000110;
    assign parity_check_matrix[426] = 10'b0100111001;
    assign parity_check_matrix[427] = 10'b1011000110;
    assign parity_check_matrix[428] = 10'b1000111001;
    assign parity_check_matrix[429] = 10'b0111000110;
    assign parity_check_matrix[430] = 10'b0011011001;
    assign parity_check_matrix[431] = 10'b1100100110;
    assign parity_check_matrix[432] = 10'b0101011001;
    assign parity_check_matrix[433] = 10'b1010100110;
    assign parity_check_matrix[434] = 10'b1001011001;
    assign parity_check_matrix[435] = 10'b0110100110;
    assign parity_check_matrix[436] = 10'b0110011001;
    assign parity_check_matrix[437] = 10'b1001100110;
    assign parity_check_matrix[438] = 10'b1010011001;
    assign parity_check_matrix[439] = 10'b0101100110;
    assign parity_check_matrix[440] = 10'b1100011001;
    assign parity_check_matrix[441] = 10'b0011100110;
    assign parity_check_matrix[442] = 10'b0011101001;
    assign parity_check_matrix[443] = 10'b1100010110;
    assign parity_check_matrix[444] = 10'b0101101001;
    assign parity_check_matrix[445] = 10'b1010010110;
    assign parity_check_matrix[446] = 10'b1001101001;
    assign parity_check_matrix[447] = 10'b0110010110;
    assign parity_check_matrix[448] = 10'b0110101001;
    assign parity_check_matrix[449] = 10'b1001010110;
    assign parity_check_matrix[450] = 10'b1010101001;
    assign parity_check_matrix[451] = 10'b0101010110;
    assign parity_check_matrix[452] = 10'b1100101001;
    assign parity_check_matrix[453] = 10'b0011010110;
    assign parity_check_matrix[454] = 10'b0111001001;
    assign parity_check_matrix[455] = 10'b1000110110;
    assign parity_check_matrix[456] = 10'b1011001001;
    assign parity_check_matrix[457] = 10'b0100110110;
    assign parity_check_matrix[458] = 10'b1101001001;
    assign parity_check_matrix[459] = 10'b0010110110;
    assign parity_check_matrix[460] = 10'b1110001001;
    assign parity_check_matrix[461] = 10'b0001110110;
    assign parity_check_matrix[462] = 10'b0011110001;
    assign parity_check_matrix[463] = 10'b1100001110;
    assign parity_check_matrix[464] = 10'b0101110001;
    assign parity_check_matrix[465] = 10'b1010001110;
    assign parity_check_matrix[466] = 10'b1001110001;
    assign parity_check_matrix[467] = 10'b0110001110;
    assign parity_check_matrix[468] = 10'b0110110001;
    assign parity_check_matrix[469] = 10'b1001001110;
    assign parity_check_matrix[470] = 10'b1010110001;
    assign parity_check_matrix[471] = 10'b0101001110;
    assign parity_check_matrix[472] = 10'b1100110001;
    assign parity_check_matrix[473] = 10'b0011001110;
    assign parity_check_matrix[474] = 10'b0111010001;
    assign parity_check_matrix[475] = 10'b1000101110;
    assign parity_check_matrix[476] = 10'b1011010001;
    assign parity_check_matrix[477] = 10'b0100101110;
    assign parity_check_matrix[478] = 10'b1101010001;
    assign parity_check_matrix[479] = 10'b0010101110;
    assign parity_check_matrix[480] = 10'b1110010001;
    assign parity_check_matrix[481] = 10'b0001101110;
    assign parity_check_matrix[482] = 10'b0111100001;
    assign parity_check_matrix[483] = 10'b1000011110;
    assign parity_check_matrix[484] = 10'b1011100001;
    assign parity_check_matrix[485] = 10'b0100011110;
    assign parity_check_matrix[486] = 10'b1101100001;
    assign parity_check_matrix[487] = 10'b0010011110;
    assign parity_check_matrix[488] = 10'b1110100001;
    assign parity_check_matrix[489] = 10'b0001011110;
    assign parity_check_matrix[490] = 10'b1111000001;
    assign parity_check_matrix[491] = 10'b0000111110;
    assign parity_check_matrix[492] = 10'b0111111111;
    assign parity_check_matrix[493] = 10'b1011111111;
    assign parity_check_matrix[494] = 10'b1101111111;
    assign parity_check_matrix[495] = 10'b1110111111;
    assign parity_check_matrix[496] = 10'b1111011111;
    assign parity_check_matrix[497] = 10'b1111101111;
    assign parity_check_matrix[498] = 10'b1111110111;
    assign parity_check_matrix[499] = 10'b1111111011;
    assign parity_check_matrix[500] = 10'b1111111101;
    assign parity_check_matrix[501] = 10'b1111111110;
    assign parity_check_matrix[502] = 10'b1000000000;
    assign parity_check_matrix[503] = 10'b0100000000;
    assign parity_check_matrix[504] = 10'b0010000000;
    assign parity_check_matrix[505] = 10'b0001000000;
    assign parity_check_matrix[506] = 10'b0000100000;
    assign parity_check_matrix[507] = 10'b0000010000;
    assign parity_check_matrix[508] = 10'b0000001000;
    assign parity_check_matrix[509] = 10'b0000000100;
    assign parity_check_matrix[510] = 10'b0000000010;
    assign parity_check_matrix[511] = 10'b0000000001;
  end else if ((CodewordWidth == 1024) && (MessageWidth == 1013)) begin : gen_1024_1013
    `BR_ASSERT_STATIC(parity_width_matches_a, ParityWidth == 11)
    assign syndrome[10] = cw[0] ^ cw[2] ^ cw[4] ^ cw[6] ^ cw[8] ^ cw[10] ^ cw[12] ^ cw[14] ^ cw[16] ^ cw[18] ^ cw[20] ^ cw[22] ^ cw[24] ^ cw[26] ^ cw[28] ^ cw[30] ^ cw[31] ^ cw[33] ^ cw[36] ^ cw[38] ^ cw[40] ^ cw[42] ^ cw[44] ^ cw[46] ^ cw[48] ^ cw[50] ^ cw[52] ^ cw[54] ^ cw[56] ^ cw[58] ^ cw[59] ^ cw[62] ^ cw[64] ^ cw[65] ^ cw[68] ^ cw[70] ^ cw[72] ^ cw[74] ^ cw[76] ^ cw[78] ^ cw[80] ^ cw[82] ^ cw[83] ^ cw[86] ^ cw[88] ^ cw[90] ^ cw[92] ^ cw[93] ^ cw[96] ^ cw[98] ^ cw[100] ^ cw[102] ^ cw[103] ^ cw[106] ^ cw[108] ^ cw[110] ^ cw[112] ^ cw[114] ^ cw[116] ^ cw[117] ^ cw[119] ^ cw[122] ^ cw[124] ^ cw[126] ^ cw[128] ^ cw[130] ^ cw[131] ^ cw[134] ^ cw[136] ^ cw[137] ^ cw[139] ^ cw[142] ^ cw[143] ^ cw[146] ^ cw[148] ^ cw[150] ^ cw[152] ^ cw[153] ^ cw[156] ^ cw[158] ^ cw[160] ^ cw[162] ^ cw[164] ^ cw[165] ^ cw[168] ^ cw[170] ^ cw[171] ^ cw[173] ^ cw[176] ^ cw[177] ^ cw[180] ^ cw[183] ^ cw[186] ^ cw[189] ^ cw[190] ^ cw[195] ^ cw[197] ^ cw[199] ^ cw[202] ^ cw[203] ^ cw[206] ^ cw[209] ^ cw[211] ^ cw[212] ^ cw[216] ^ cw[217] ^ cw[222] ^ cw[225] ^ cw[227] ^ cw[229] ^ cw[232] ^ cw[233] ^ cw[235] ^ cw[237] ^ cw[241] ^ cw[244] ^ cw[246] ^ cw[248] ^ cw[252] ^ cw[253] ^ cw[256] ^ cw[260] ^ cw[262] ^ cw[263] ^ cw[268] ^ cw[270] ^ cw[272] ^ cw[276] ^ cw[278] ^ cw[281] ^ cw[282] ^ cw[285] ^ cw[288] ^ cw[290] ^ cw[294] ^ cw[295] ^ cw[296] ^ cw[299] ^ cw[302] ^ cw[303] ^ cw[306] ^ cw[308] ^ cw[311] ^ cw[313] ^ cw[315] ^ cw[317] ^ cw[319] ^ cw[321] ^ cw[323] ^ cw[325] ^ cw[326] ^ cw[329] ^ cw[331] ^ cw[332] ^ cw[335] ^ cw[337] ^ cw[339] ^ cw[341] ^ cw[343] ^ cw[345] ^ cw[346] ^ cw[349] ^ cw[351] ^ cw[352] ^ cw[355] ^ cw[357] ^ cw[359] ^ cw[361] ^ cw[362] ^ cw[365] ^ cw[367] ^ cw[368] ^ cw[371] ^ cw[373] ^ cw[374] ^ cw[377] ^ cw[379] ^ cw[380] ^ cw[382] ^ cw[385] ^ cw[386] ^ cw[388] ^ cw[391] ^ cw[392] ^ cw[395] ^ cw[397] ^ cw[399] ^ cw[401] ^ cw[403] ^ cw[405] ^ cw[407] ^ cw[409] ^ cw[410] ^ cw[412] ^ cw[415] ^ cw[417] ^ cw[419] ^ cw[421] ^ cw[423] ^ cw[425] ^ cw[427] ^ cw[428] ^ cw[431] ^ cw[433] ^ cw[434] ^ cw[437] ^ cw[439] ^ cw[440] ^ cw[442] ^ cw[445] ^ cw[447] ^ cw[448] ^ cw[450] ^ cw[452] ^ cw[454] ^ cw[457] ^ cw[459] ^ cw[461] ^ cw[463] ^ cw[465] ^ cw[467] ^ cw[468] ^ cw[471] ^ cw[473] ^ cw[475] ^ cw[477] ^ cw[478] ^ cw[480] ^ cw[483] ^ cw[485] ^ cw[486] ^ cw[488] ^ cw[491] ^ cw[492] ^ cw[494] ^ cw[497] ^ cw[499] ^ cw[501] ^ cw[503] ^ cw[504] ^ cw[507] ^ cw[509] ^ cw[510] ^ cw[512] ^ cw[515] ^ cw[516] ^ cw[519] ^ cw[521] ^ cw[523] ^ cw[524] ^ cw[526] ^ cw[528] ^ cw[530] ^ cw[532] ^ cw[535] ^ cw[537] ^ cw[539] ^ cw[541] ^ cw[542] ^ cw[545] ^ cw[547] ^ cw[549] ^ cw[550] ^ cw[552] ^ cw[554] ^ cw[557] ^ cw[558] ^ cw[560] ^ cw[562] ^ cw[564] ^ cw[566] ^ cw[568] ^ cw[570] ^ cw[572] ^ cw[574] ^ cw[575] ^ cw[578] ^ cw[580] ^ cw[581] ^ cw[584] ^ cw[586] ^ cw[588] ^ cw[590] ^ cw[592] ^ cw[593] ^ cw[595] ^ cw[598] ^ cw[600] ^ cw[601] ^ cw[604] ^ cw[605] ^ cw[608] ^ cw[610] ^ cw[611] ^ cw[614] ^ cw[616] ^ cw[618] ^ cw[620] ^ cw[622] ^ cw[623] ^ cw[625] ^ cw[628] ^ cw[630] ^ cw[631] ^ cw[633] ^ cw[635] ^ cw[638] ^ cw[640] ^ cw[642] ^ cw[644] ^ cw[645] ^ cw[648] ^ cw[650] ^ cw[652] ^ cw[653] ^ cw[655] ^ cw[658] ^ cw[660] ^ cw[661] ^ cw[664] ^ cw[666] ^ cw[668] ^ cw[670] ^ cw[671] ^ cw[673] ^ cw[676] ^ cw[678] ^ cw[680] ^ cw[681] ^ cw[683] ^ cw[685] ^ cw[688] ^ cw[690] ^ cw[691] ^ cw[693] ^ cw[695] ^ cw[697] ^ cw[700] ^ cw[702] ^ cw[704] ^ cw[705] ^ cw[708] ^ cw[710] ^ cw[711] ^ cw[714] ^ cw[716] ^ cw[718] ^ cw[720] ^ cw[721] ^ cw[723] ^ cw[726] ^ cw[728] ^ cw[730] ^ cw[731] ^ cw[733] ^ cw[735] ^ cw[738] ^ cw[740] ^ cw[741] ^ cw[744] ^ cw[745] ^ cw[747] ^ cw[750] ^ cw[752] ^ cw[754] ^ cw[755] ^ cw[757] ^ cw[759] ^ cw[762] ^ cw[764] ^ cw[765] ^ cw[767] ^ cw[769] ^ cw[771] ^ cw[774] ^ cw[775] ^ cw[777] ^ cw[780] ^ cw[781] ^ cw[783] ^ cw[785] ^ cw[788] ^ cw[790] ^ cw[792] ^ cw[794] ^ cw[795] ^ cw[797] ^ cw[800] ^ cw[802] ^ cw[803] ^ cw[805] ^ cw[807] ^ cw[809] ^ cw[812] ^ cw[814] ^ cw[816] ^ cw[818] ^ cw[819] ^ cw[821] ^ cw[822] ^ cw[825] ^ cw[827] ^ cw[829] ^ cw[830] ^ cw[832] ^ cw[834] ^ cw[836] ^ cw[837] ^ cw[839] ^ cw[841] ^ cw[843] ^ cw[845] ^ cw[846] ^ cw[847] ^ cw[849] ^ cw[852] ^ cw[853] ^ cw[855] ^ cw[856] ^ cw[859] ^ cw[860] ^ cw[862] ^ cw[864] ^ cw[865] ^ cw[866] ^ cw[869] ^ cw[870] ^ cw[872] ^ cw[875] ^ cw[877] ^ cw[878] ^ cw[880] ^ cw[881] ^ cw[882] ^ cw[884] ^ cw[886] ^ cw[887] ^ cw[889] ^ cw[892] ^ cw[893] ^ cw[895] ^ cw[896] ^ cw[898] ^ cw[899] ^ cw[901] ^ cw[902] ^ cw[906] ^ cw[907] ^ cw[908] ^ cw[911] ^ cw[912] ^ cw[915] ^ cw[916] ^ cw[917] ^ cw[919] ^ cw[922] ^ cw[924] ^ cw[926] ^ cw[927] ^ cw[928] ^ cw[931] ^ cw[933] ^ cw[934] ^ cw[936] ^ cw[938] ^ cw[940] ^ cw[942] ^ cw[943] ^ cw[945] ^ cw[947] ^ cw[948] ^ cw[950] ^ cw[951] ^ cw[953] ^ cw[955] ^ cw[957] ^ cw[958] ^ cw[960] ^ cw[963] ^ cw[964] ^ cw[966] ^ cw[967] ^ cw[968] ^ cw[970] ^ cw[972] ^ cw[973] ^ cw[975] ^ cw[976] ^ cw[978] ^ cw[979] ^ cw[982] ^ cw[983] ^ cw[984] ^ cw[986] ^ cw[988] ^ cw[990] ^ cw[991] ^ cw[993] ^ cw[995] ^ cw[996] ^ cw[997] ^ cw[1000] ^ cw[1001] ^ cw[1002] ^ cw[1004] ^ cw[1005] ^ cw[1006] ^ cw[1008] ^ cw[1009] ^ cw[1011] ^ cw[1012] ^ cw[1013];
    assign syndrome[9] = cw[0] ^ cw[2] ^ cw[4] ^ cw[6] ^ cw[8] ^ cw[10] ^ cw[12] ^ cw[14] ^ cw[16] ^ cw[18] ^ cw[20] ^ cw[22] ^ cw[24] ^ cw[26] ^ cw[27] ^ cw[29] ^ cw[32] ^ cw[34] ^ cw[36] ^ cw[38] ^ cw[40] ^ cw[42] ^ cw[44] ^ cw[46] ^ cw[48] ^ cw[50] ^ cw[52] ^ cw[54] ^ cw[55] ^ cw[58] ^ cw[60] ^ cw[61] ^ cw[64] ^ cw[66] ^ cw[68] ^ cw[70] ^ cw[72] ^ cw[74] ^ cw[76] ^ cw[78] ^ cw[79] ^ cw[82] ^ cw[84] ^ cw[86] ^ cw[88] ^ cw[89] ^ cw[92] ^ cw[94] ^ cw[96] ^ cw[98] ^ cw[99] ^ cw[102] ^ cw[104] ^ cw[106] ^ cw[108] ^ cw[110] ^ cw[112] ^ cw[113] ^ cw[115] ^ cw[118] ^ cw[120] ^ cw[122] ^ cw[124] ^ cw[126] ^ cw[127] ^ cw[130] ^ cw[132] ^ cw[133] ^ cw[135] ^ cw[138] ^ cw[140] ^ cw[142] ^ cw[143] ^ cw[146] ^ cw[148] ^ cw[149] ^ cw[152] ^ cw[154] ^ cw[156] ^ cw[158] ^ cw[160] ^ cw[161] ^ cw[164] ^ cw[166] ^ cw[167] ^ cw[169] ^ cw[172] ^ cw[174] ^ cw[176] ^ cw[177] ^ cw[180] ^ cw[183] ^ cw[186] ^ cw[187] ^ cw[191] ^ cw[195] ^ cw[197] ^ cw[199] ^ cw[202] ^ cw[204] ^ cw[206] ^ cw[208] ^ cw[211] ^ cw[213] ^ cw[214] ^ cw[219] ^ cw[221] ^ cw[224] ^ cw[227] ^ cw[228] ^ cw[230] ^ cw[234] ^ cw[236] ^ cw[238] ^ cw[241] ^ cw[243] ^ cw[247] ^ cw[249] ^ cw[250] ^ cw[254] ^ cw[256] ^ cw[260] ^ cw[262] ^ cw[265] ^ cw[267] ^ cw[269] ^ cw[273] ^ cw[275] ^ cw[279] ^ cw[280] ^ cw[283] ^ cw[285] ^ cw[288] ^ cw[291] ^ cw[292] ^ cw[295] ^ cw[298] ^ cw[299] ^ cw[301] ^ cw[305] ^ cw[306] ^ cw[308] ^ cw[311] ^ cw[313] ^ cw[315] ^ cw[317] ^ cw[319] ^ cw[321] ^ cw[322] ^ cw[325] ^ cw[327] ^ cw[328] ^ cw[331] ^ cw[333] ^ cw[335] ^ cw[337] ^ cw[339] ^ cw[341] ^ cw[342] ^ cw[345] ^ cw[347] ^ cw[348] ^ cw[351] ^ cw[353] ^ cw[355] ^ cw[357] ^ cw[358] ^ cw[361] ^ cw[363] ^ cw[364] ^ cw[367] ^ cw[369] ^ cw[370] ^ cw[373] ^ cw[375] ^ cw[376] ^ cw[378] ^ cw[381] ^ cw[383] ^ cw[384] ^ cw[386] ^ cw[389] ^ cw[391] ^ cw[392] ^ cw[395] ^ cw[397] ^ cw[399] ^ cw[401] ^ cw[403] ^ cw[405] ^ cw[406] ^ cw[408] ^ cw[411] ^ cw[413] ^ cw[415] ^ cw[417] ^ cw[419] ^ cw[421] ^ cw[422] ^ cw[424] ^ cw[427] ^ cw[429] ^ cw[431] ^ cw[433] ^ cw[435] ^ cw[436] ^ cw[438] ^ cw[441] ^ cw[443] ^ cw[444] ^ cw[446] ^ cw[449] ^ cw[451] ^ cw[452] ^ cw[454] ^ cw[457] ^ cw[459] ^ cw[461] ^ cw[463] ^ cw[464] ^ cw[467] ^ cw[469] ^ cw[471] ^ cw[473] ^ cw[474] ^ cw[476] ^ cw[479] ^ cw[481] ^ cw[483] ^ cw[484] ^ cw[487] ^ cw[489] ^ cw[490] ^ cw[492] ^ cw[494] ^ cw[497] ^ cw[499] ^ cw[500] ^ cw[503] ^ cw[505] ^ cw[506] ^ cw[508] ^ cw[511] ^ cw[513] ^ cw[515] ^ cw[516] ^ cw[518] ^ cw[520] ^ cw[522] ^ cw[525] ^ cw[527] ^ cw[528] ^ cw[530] ^ cw[532] ^ cw[534] ^ cw[537] ^ cw[538] ^ cw[541] ^ cw[543] ^ cw[545] ^ cw[546] ^ cw[548] ^ cw[551] ^ cw[553] ^ cw[554] ^ cw[557] ^ cw[558] ^ cw[560] ^ cw[562] ^ cw[564] ^ cw[566] ^ cw[568] ^ cw[570] ^ cw[571] ^ cw[573] ^ cw[576] ^ cw[578] ^ cw[580] ^ cw[582] ^ cw[584] ^ cw[586] ^ cw[588] ^ cw[589] ^ cw[591] ^ cw[594] ^ cw[596] ^ cw[597] ^ cw[600] ^ cw[602] ^ cw[604] ^ cw[605] ^ cw[607] ^ cw[610] ^ cw[612] ^ cw[613] ^ cw[616] ^ cw[618] ^ cw[619] ^ cw[622] ^ cw[624] ^ cw[626] ^ cw[627] ^ cw[629] ^ cw[632] ^ cw[634] ^ cw[635] ^ cw[638] ^ cw[640] ^ cw[641] ^ cw[644] ^ cw[646] ^ cw[648] ^ cw[649] ^ cw[651] ^ cw[654] ^ cw[656] ^ cw[658] ^ cw[660] ^ cw[661] ^ cw[664] ^ cw[666] ^ cw[667] ^ cw[669] ^ cw[672] ^ cw[674] ^ cw[676] ^ cw[677] ^ cw[679] ^ cw[682] ^ cw[684] ^ cw[685] ^ cw[687] ^ cw[689] ^ cw[692] ^ cw[694] ^ cw[695] ^ cw[697] ^ cw[700] ^ cw[702] ^ cw[704] ^ cw[705] ^ cw[707] ^ cw[710] ^ cw[712] ^ cw[714] ^ cw[716] ^ cw[717] ^ cw[719] ^ cw[722] ^ cw[724] ^ cw[726] ^ cw[727] ^ cw[729] ^ cw[732] ^ cw[734] ^ cw[735] ^ cw[737] ^ cw[740] ^ cw[742] ^ cw[743] ^ cw[745] ^ cw[748] ^ cw[750] ^ cw[751] ^ cw[753] ^ cw[756] ^ cw[758] ^ cw[759] ^ cw[761] ^ cw[763] ^ cw[766] ^ cw[768] ^ cw[769] ^ cw[771] ^ cw[773] ^ cw[775] ^ cw[778] ^ cw[779] ^ cw[781] ^ cw[784] ^ cw[785] ^ cw[788] ^ cw[790] ^ cw[791] ^ cw[793] ^ cw[796] ^ cw[798] ^ cw[799] ^ cw[801] ^ cw[804] ^ cw[806] ^ cw[807] ^ cw[809] ^ cw[812] ^ cw[814] ^ cw[815] ^ cw[818] ^ cw[819] ^ cw[821] ^ cw[823] ^ cw[824] ^ cw[827] ^ cw[829] ^ cw[830] ^ cw[831] ^ cw[834] ^ cw[835] ^ cw[837] ^ cw[839] ^ cw[841] ^ cw[842] ^ cw[844] ^ cw[847] ^ cw[848] ^ cw[850] ^ cw[851] ^ cw[854] ^ cw[855] ^ cw[857] ^ cw[859] ^ cw[861] ^ cw[862] ^ cw[863] ^ cw[865] ^ cw[867] ^ cw[869] ^ cw[871] ^ cw[872] ^ cw[874] ^ cw[877] ^ cw[878] ^ cw[879] ^ cw[881] ^ cw[883] ^ cw[884] ^ cw[885] ^ cw[887] ^ cw[889] ^ cw[891] ^ cw[893] ^ cw[894] ^ cw[896] ^ cw[897] ^ cw[899] ^ cw[902] ^ cw[903] ^ cw[905] ^ cw[907] ^ cw[909] ^ cw[911] ^ cw[913] ^ cw[914] ^ cw[915] ^ cw[917] ^ cw[919] ^ cw[920] ^ cw[924] ^ cw[925] ^ cw[927] ^ cw[929] ^ cw[931] ^ cw[932] ^ cw[934] ^ cw[935] ^ cw[937] ^ cw[940] ^ cw[941] ^ cw[942] ^ cw[944] ^ cw[946] ^ cw[948] ^ cw[950] ^ cw[952] ^ cw[954] ^ cw[955] ^ cw[956] ^ cw[958] ^ cw[959] ^ cw[960] ^ cw[962] ^ cw[966] ^ cw[967] ^ cw[969] ^ cw[970] ^ cw[971] ^ cw[973] ^ cw[975] ^ cw[977] ^ cw[978] ^ cw[979] ^ cw[982] ^ cw[983] ^ cw[985] ^ cw[987] ^ cw[988] ^ cw[989] ^ cw[992] ^ cw[993] ^ cw[994] ^ cw[996] ^ cw[998] ^ cw[999] ^ cw[1001] ^ cw[1002] ^ cw[1003] ^ cw[1005] ^ cw[1007] ^ cw[1008] ^ cw[1009] ^ cw[1010] ^ cw[1012] ^ cw[1014];
    assign syndrome[8] = cw[0] ^ cw[2] ^ cw[4] ^ cw[6] ^ cw[8] ^ cw[10] ^ cw[12] ^ cw[14] ^ cw[16] ^ cw[18] ^ cw[20] ^ cw[22] ^ cw[23] ^ cw[25] ^ cw[28] ^ cw[30] ^ cw[32] ^ cw[34] ^ cw[36] ^ cw[38] ^ cw[40] ^ cw[42] ^ cw[44] ^ cw[46] ^ cw[48] ^ cw[50] ^ cw[51] ^ cw[54] ^ cw[56] ^ cw[57] ^ cw[60] ^ cw[62] ^ cw[64] ^ cw[66] ^ cw[68] ^ cw[70] ^ cw[72] ^ cw[74] ^ cw[75] ^ cw[78] ^ cw[80] ^ cw[82] ^ cw[84] ^ cw[85] ^ cw[88] ^ cw[90] ^ cw[92] ^ cw[94] ^ cw[95] ^ cw[98] ^ cw[100] ^ cw[102] ^ cw[104] ^ cw[106] ^ cw[108] ^ cw[109] ^ cw[111] ^ cw[114] ^ cw[116] ^ cw[118] ^ cw[120] ^ cw[122] ^ cw[123] ^ cw[126] ^ cw[128] ^ cw[129] ^ cw[132] ^ cw[134] ^ cw[135] ^ cw[138] ^ cw[139] ^ cw[142] ^ cw[144] ^ cw[145] ^ cw[148] ^ cw[150] ^ cw[152] ^ cw[154] ^ cw[156] ^ cw[157] ^ cw[160] ^ cw[162] ^ cw[163] ^ cw[166] ^ cw[168] ^ cw[169] ^ cw[172] ^ cw[173] ^ cw[176] ^ cw[178] ^ cw[180] ^ cw[183] ^ cw[184] ^ cw[188] ^ cw[192] ^ cw[195] ^ cw[197] ^ cw[199] ^ cw[202] ^ cw[204] ^ cw[205] ^ cw[207] ^ cw[211] ^ cw[213] ^ cw[216] ^ cw[218] ^ cw[221] ^ cw[223] ^ cw[226] ^ cw[229] ^ cw[231] ^ cw[234] ^ cw[236] ^ cw[239] ^ cw[240] ^ cw[244] ^ cw[247] ^ cw[249] ^ cw[250] ^ cw[253] ^ cw[257] ^ cw[260] ^ cw[261] ^ cw[264] ^ cw[266] ^ cw[271] ^ cw[273] ^ cw[275] ^ cw[278] ^ cw[281] ^ cw[282] ^ cw[286] ^ cw[287] ^ cw[291] ^ cw[292] ^ cw[295] ^ cw[296] ^ cw[300] ^ cw[301] ^ cw[303] ^ cw[307] ^ cw[308] ^ cw[311] ^ cw[313] ^ cw[315] ^ cw[317] ^ cw[318] ^ cw[321] ^ cw[323] ^ cw[324] ^ cw[327] ^ cw[329] ^ cw[331] ^ cw[333] ^ cw[335] ^ cw[337] ^ cw[338] ^ cw[341] ^ cw[343] ^ cw[344] ^ cw[347] ^ cw[349] ^ cw[351] ^ cw[353] ^ cw[354] ^ cw[357] ^ cw[359] ^ cw[360] ^ cw[363] ^ cw[365] ^ cw[366] ^ cw[369] ^ cw[371] ^ cw[372] ^ cw[375] ^ cw[377] ^ cw[378] ^ cw[381] ^ cw[382] ^ cw[384] ^ cw[387] ^ cw[388] ^ cw[391] ^ cw[393] ^ cw[395] ^ cw[397] ^ cw[399] ^ cw[401] ^ cw[402] ^ cw[404] ^ cw[407] ^ cw[409] ^ cw[411] ^ cw[413] ^ cw[415] ^ cw[417] ^ cw[418] ^ cw[420] ^ cw[423] ^ cw[425] ^ cw[427] ^ cw[429] ^ cw[430] ^ cw[432] ^ cw[435] ^ cw[437] ^ cw[439] ^ cw[441] ^ cw[443] ^ cw[444] ^ cw[446] ^ cw[448] ^ cw[450] ^ cw[453] ^ cw[455] ^ cw[457] ^ cw[459] ^ cw[460] ^ cw[462] ^ cw[465] ^ cw[467] ^ cw[469] ^ cw[470] ^ cw[472] ^ cw[475] ^ cw[477] ^ cw[479] ^ cw[481] ^ cw[482] ^ cw[484] ^ cw[487] ^ cw[488] ^ cw[490] ^ cw[493] ^ cw[495] ^ cw[496] ^ cw[499] ^ cw[501] ^ cw[502] ^ cw[505] ^ cw[507] ^ cw[508] ^ cw[511] ^ cw[512] ^ cw[514] ^ cw[517] ^ cw[519] ^ cw[520] ^ cw[522] ^ cw[524] ^ cw[526] ^ cw[529] ^ cw[531] ^ cw[532] ^ cw[535] ^ cw[537] ^ cw[538] ^ cw[541] ^ cw[542] ^ cw[544] ^ cw[546] ^ cw[549] ^ cw[550] ^ cw[553] ^ cw[555] ^ cw[557] ^ cw[558] ^ cw[560] ^ cw[562] ^ cw[564] ^ cw[565] ^ cw[567] ^ cw[570] ^ cw[572] ^ cw[574] ^ cw[576] ^ cw[578] ^ cw[580] ^ cw[582] ^ cw[584] ^ cw[585] ^ cw[587] ^ cw[590] ^ cw[592] ^ cw[594] ^ cw[596] ^ cw[597] ^ cw[600] ^ cw[601] ^ cw[603] ^ cw[606] ^ cw[608] ^ cw[609] ^ cw[612] ^ cw[614] ^ cw[615] ^ cw[618] ^ cw[620] ^ cw[621] ^ cw[624] ^ cw[626] ^ cw[627] ^ cw[630] ^ cw[631] ^ cw[634] ^ cw[636] ^ cw[637] ^ cw[640] ^ cw[642] ^ cw[644] ^ cw[646] ^ cw[647] ^ cw[649] ^ cw[652] ^ cw[653] ^ cw[656] ^ cw[658] ^ cw[660] ^ cw[662] ^ cw[663] ^ cw[665] ^ cw[668] ^ cw[670] ^ cw[672] ^ cw[674] ^ cw[675] ^ cw[677] ^ cw[680] ^ cw[681] ^ cw[684] ^ cw[686] ^ cw[687] ^ cw[689] ^ cw[691] ^ cw[693] ^ cw[696] ^ cw[698] ^ cw[700] ^ cw[701] ^ cw[703] ^ cw[705] ^ cw[708] ^ cw[710] ^ cw[712] ^ cw[713] ^ cw[715] ^ cw[718] ^ cw[720] ^ cw[722] ^ cw[724] ^ cw[725] ^ cw[727] ^ cw[730] ^ cw[731] ^ cw[734] ^ cw[736] ^ cw[737] ^ cw[739] ^ cw[741] ^ cw[744] ^ cw[746] ^ cw[748] ^ cw[749] ^ cw[751] ^ cw[754] ^ cw[755] ^ cw[758] ^ cw[760] ^ cw[761] ^ cw[763] ^ cw[765] ^ cw[767] ^ cw[770] ^ cw[772] ^ cw[773] ^ cw[775] ^ cw[777] ^ cw[780] ^ cw[782] ^ cw[784] ^ cw[785] ^ cw[787] ^ cw[789] ^ cw[792] ^ cw[794] ^ cw[796] ^ cw[798] ^ cw[799] ^ cw[801] ^ cw[803] ^ cw[805] ^ cw[808] ^ cw[810] ^ cw[812] ^ cw[813] ^ cw[815] ^ cw[818] ^ cw[819] ^ cw[820] ^ cw[822] ^ cw[825] ^ cw[827] ^ cw[828] ^ cw[830] ^ cw[832] ^ cw[833] ^ cw[835] ^ cw[837] ^ cw[838] ^ cw[841] ^ cw[843] ^ cw[845] ^ cw[847] ^ cw[848] ^ cw[850] ^ cw[852] ^ cw[853] ^ cw[854] ^ cw[857] ^ cw[858] ^ cw[861] ^ cw[862] ^ cw[864] ^ cw[865] ^ cw[866] ^ cw[868] ^ cw[871] ^ cw[873] ^ cw[875] ^ cw[876] ^ cw[878] ^ cw[879] ^ cw[880] ^ cw[882] ^ cw[885] ^ cw[886] ^ cw[888] ^ cw[890] ^ cw[891] ^ cw[892] ^ cw[894] ^ cw[896] ^ cw[898] ^ cw[899] ^ cw[902] ^ cw[903] ^ cw[904] ^ cw[907] ^ cw[908] ^ cw[911] ^ cw[912] ^ cw[914] ^ cw[916] ^ cw[918] ^ cw[919] ^ cw[921] ^ cw[923] ^ cw[926] ^ cw[927] ^ cw[929] ^ cw[930] ^ cw[932] ^ cw[933] ^ cw[935] ^ cw[938] ^ cw[939] ^ cw[941] ^ cw[942] ^ cw[944] ^ cw[947] ^ cw[949] ^ cw[950] ^ cw[952] ^ cw[953] ^ cw[956] ^ cw[957] ^ cw[958] ^ cw[959] ^ cw[960] ^ cw[963] ^ cw[965] ^ cw[967] ^ cw[968] ^ cw[970] ^ cw[972] ^ cw[973] ^ cw[974] ^ cw[977] ^ cw[978] ^ cw[980] ^ cw[981] ^ cw[982] ^ cw[985] ^ cw[986] ^ cw[989] ^ cw[990] ^ cw[992] ^ cw[994] ^ cw[995] ^ cw[997] ^ cw[998] ^ cw[999] ^ cw[1000] ^ cw[1002] ^ cw[1004] ^ cw[1005] ^ cw[1006] ^ cw[1007] ^ cw[1009] ^ cw[1010] ^ cw[1011] ^ cw[1015];
    assign syndrome[7] = cw[0] ^ cw[2] ^ cw[4] ^ cw[6] ^ cw[8] ^ cw[10] ^ cw[12] ^ cw[14] ^ cw[16] ^ cw[18] ^ cw[19] ^ cw[21] ^ cw[24] ^ cw[26] ^ cw[28] ^ cw[30] ^ cw[32] ^ cw[34] ^ cw[36] ^ cw[38] ^ cw[40] ^ cw[42] ^ cw[44] ^ cw[46] ^ cw[47] ^ cw[50] ^ cw[52] ^ cw[53] ^ cw[56] ^ cw[58] ^ cw[60] ^ cw[62] ^ cw[64] ^ cw[66] ^ cw[68] ^ cw[70] ^ cw[71] ^ cw[74] ^ cw[76] ^ cw[78] ^ cw[80] ^ cw[81] ^ cw[84] ^ cw[86] ^ cw[88] ^ cw[90] ^ cw[91] ^ cw[94] ^ cw[96] ^ cw[98] ^ cw[100] ^ cw[102] ^ cw[104] ^ cw[105] ^ cw[107] ^ cw[110] ^ cw[112] ^ cw[114] ^ cw[116] ^ cw[118] ^ cw[120] ^ cw[122] ^ cw[123] ^ cw[125] ^ cw[127] ^ cw[130] ^ cw[131] ^ cw[134] ^ cw[136] ^ cw[138] ^ cw[140] ^ cw[141] ^ cw[144] ^ cw[146] ^ cw[148] ^ cw[150] ^ cw[152] ^ cw[154] ^ cw[156] ^ cw[157] ^ cw[159] ^ cw[161] ^ cw[164] ^ cw[165] ^ cw[168] ^ cw[170] ^ cw[172] ^ cw[174] ^ cw[176] ^ cw[178] ^ cw[180] ^ cw[181] ^ cw[185] ^ cw[189] ^ cw[192] ^ cw[194] ^ cw[197] ^ cw[199] ^ cw[200] ^ cw[204] ^ cw[206] ^ cw[209] ^ cw[210] ^ cw[213] ^ cw[215] ^ cw[219] ^ cw[220] ^ cw[224] ^ cw[227] ^ cw[229] ^ cw[231] ^ cw[233] ^ cw[236] ^ cw[239] ^ cw[240] ^ cw[243] ^ cw[247] ^ cw[248] ^ cw[251] ^ cw[255] ^ cw[258] ^ cw[259] ^ cw[262] ^ cw[264] ^ cw[266] ^ cw[269] ^ cw[272] ^ cw[276] ^ cw[277] ^ cw[280] ^ cw[283] ^ cw[286] ^ cw[289] ^ cw[290] ^ cw[294] ^ cw[295] ^ cw[297] ^ cw[300] ^ cw[301] ^ cw[303] ^ cw[306] ^ cw[309] ^ cw[311] ^ cw[313] ^ cw[314] ^ cw[317] ^ cw[319] ^ cw[320] ^ cw[323] ^ cw[325] ^ cw[327] ^ cw[329] ^ cw[331] ^ cw[333] ^ cw[334] ^ cw[337] ^ cw[339] ^ cw[340] ^ cw[343] ^ cw[345] ^ cw[347] ^ cw[349] ^ cw[350] ^ cw[353] ^ cw[355] ^ cw[356] ^ cw[359] ^ cw[361] ^ cw[363] ^ cw[365] ^ cw[366] ^ cw[369] ^ cw[370] ^ cw[372] ^ cw[374] ^ cw[376] ^ cw[379] ^ cw[380] ^ cw[383] ^ cw[385] ^ cw[387] ^ cw[389] ^ cw[391] ^ cw[393] ^ cw[395] ^ cw[397] ^ cw[398] ^ cw[400] ^ cw[403] ^ cw[405] ^ cw[407] ^ cw[409] ^ cw[411] ^ cw[413] ^ cw[415] ^ cw[416] ^ cw[419] ^ cw[421] ^ cw[423] ^ cw[425] ^ cw[426] ^ cw[429] ^ cw[431] ^ cw[432] ^ cw[435] ^ cw[436] ^ cw[438] ^ cw[440] ^ cw[442] ^ cw[445] ^ cw[447] ^ cw[449] ^ cw[451] ^ cw[453] ^ cw[455] ^ cw[456] ^ cw[458] ^ cw[461] ^ cw[463] ^ cw[465] ^ cw[466] ^ cw[469] ^ cw[471] ^ cw[472] ^ cw[475] ^ cw[476] ^ cw[479] ^ cw[480] ^ cw[482] ^ cw[485] ^ cw[486] ^ cw[489] ^ cw[491] ^ cw[493] ^ cw[495] ^ cw[496] ^ cw[498] ^ cw[500] ^ cw[503] ^ cw[504] ^ cw[507] ^ cw[509] ^ cw[511] ^ cw[513] ^ cw[514] ^ cw[517] ^ cw[518] ^ cw[520] ^ cw[523] ^ cw[524] ^ cw[527] ^ cw[528] ^ cw[531] ^ cw[533] ^ cw[534] ^ cw[537] ^ cw[539] ^ cw[540] ^ cw[543] ^ cw[545] ^ cw[546] ^ cw[549] ^ cw[550] ^ cw[553] ^ cw[554] ^ cw[557] ^ cw[558] ^ cw[560] ^ cw[561] ^ cw[563] ^ cw[566] ^ cw[568] ^ cw[570] ^ cw[572] ^ cw[574] ^ cw[576] ^ cw[577] ^ cw[580] ^ cw[582] ^ cw[583] ^ cw[585] ^ cw[588] ^ cw[589] ^ cw[592] ^ cw[593] ^ cw[596] ^ cw[598] ^ cw[599] ^ cw[602] ^ cw[604] ^ cw[606] ^ cw[608] ^ cw[610] ^ cw[612] ^ cw[614] ^ cw[615] ^ cw[617] ^ cw[619] ^ cw[622] ^ cw[623] ^ cw[626] ^ cw[628] ^ cw[630] ^ cw[632] ^ cw[634] ^ cw[636] ^ cw[637] ^ cw[640] ^ cw[641] ^ cw[643] ^ cw[645] ^ cw[648] ^ cw[650] ^ cw[652] ^ cw[654] ^ cw[656] ^ cw[657] ^ cw[659] ^ cw[662] ^ cw[664] ^ cw[665] ^ cw[668] ^ cw[669] ^ cw[672] ^ cw[673] ^ cw[675] ^ cw[678] ^ cw[679] ^ cw[682] ^ cw[683] ^ cw[686] ^ cw[688] ^ cw[689] ^ cw[692] ^ cw[693] ^ cw[696] ^ cw[697] ^ cw[699] ^ cw[702] ^ cw[704] ^ cw[706] ^ cw[708] ^ cw[709] ^ cw[712] ^ cw[714] ^ cw[715] ^ cw[718] ^ cw[719] ^ cw[722] ^ cw[723] ^ cw[725] ^ cw[728] ^ cw[729] ^ cw[732] ^ cw[733] ^ cw[736] ^ cw[738] ^ cw[739] ^ cw[742] ^ cw[743] ^ cw[746] ^ cw[747] ^ cw[749] ^ cw[752] ^ cw[753] ^ cw[756] ^ cw[757] ^ cw[760] ^ cw[762] ^ cw[763] ^ cw[766] ^ cw[767] ^ cw[770] ^ cw[771] ^ cw[773] ^ cw[776] ^ cw[777] ^ cw[780] ^ cw[781] ^ cw[784] ^ cw[786] ^ cw[787] ^ cw[789] ^ cw[791] ^ cw[793] ^ cw[795] ^ cw[797] ^ cw[800] ^ cw[802] ^ cw[804] ^ cw[806] ^ cw[808] ^ cw[810] ^ cw[811] ^ cw[813] ^ cw[815] ^ cw[817] ^ cw[819] ^ cw[821] ^ cw[822] ^ cw[825] ^ cw[827] ^ cw[829] ^ cw[830] ^ cw[831] ^ cw[833] ^ cw[835] ^ cw[837] ^ cw[838] ^ cw[840] ^ cw[843] ^ cw[844] ^ cw[846] ^ cw[848] ^ cw[850] ^ cw[851] ^ cw[853] ^ cw[855] ^ cw[856] ^ cw[858] ^ cw[860] ^ cw[862] ^ cw[863] ^ cw[865] ^ cw[867] ^ cw[869] ^ cw[870] ^ cw[873] ^ cw[875] ^ cw[876] ^ cw[877] ^ cw[880] ^ cw[881] ^ cw[883] ^ cw[885] ^ cw[886] ^ cw[888] ^ cw[889] ^ cw[890] ^ cw[892] ^ cw[893] ^ cw[896] ^ cw[897] ^ cw[900] ^ cw[902] ^ cw[903] ^ cw[905] ^ cw[906] ^ cw[909] ^ cw[910] ^ cw[912] ^ cw[914] ^ cw[916] ^ cw[917] ^ cw[918] ^ cw[922] ^ cw[923] ^ cw[925] ^ cw[927] ^ cw[928] ^ cw[930] ^ cw[932] ^ cw[934] ^ cw[936] ^ cw[938] ^ cw[939] ^ cw[940] ^ cw[943] ^ cw[944] ^ cw[946] ^ cw[947] ^ cw[949] ^ cw[951] ^ cw[952] ^ cw[954] ^ cw[955] ^ cw[959] ^ cw[960] ^ cw[961] ^ cw[962] ^ cw[964] ^ cw[967] ^ cw[968] ^ cw[970] ^ cw[971] ^ cw[972] ^ cw[974] ^ cw[976] ^ cw[978] ^ cw[980] ^ cw[982] ^ cw[983] ^ cw[984] ^ cw[987] ^ cw[989] ^ cw[990] ^ cw[991] ^ cw[994] ^ cw[995] ^ cw[997] ^ cw[998] ^ cw[999] ^ cw[1000] ^ cw[1001] ^ cw[1003] ^ cw[1004] ^ cw[1007] ^ cw[1008] ^ cw[1010] ^ cw[1011] ^ cw[1012] ^ cw[1016];
    assign syndrome[6] = cw[0] ^ cw[2] ^ cw[4] ^ cw[6] ^ cw[8] ^ cw[10] ^ cw[12] ^ cw[14] ^ cw[15] ^ cw[17] ^ cw[20] ^ cw[22] ^ cw[24] ^ cw[26] ^ cw[28] ^ cw[30] ^ cw[32] ^ cw[34] ^ cw[36] ^ cw[38] ^ cw[40] ^ cw[42] ^ cw[43] ^ cw[46] ^ cw[48] ^ cw[49] ^ cw[52] ^ cw[54] ^ cw[56] ^ cw[58] ^ cw[60] ^ cw[62] ^ cw[64] ^ cw[66] ^ cw[67] ^ cw[70] ^ cw[72] ^ cw[74] ^ cw[76] ^ cw[77] ^ cw[80] ^ cw[82] ^ cw[84] ^ cw[86] ^ cw[87] ^ cw[90] ^ cw[92] ^ cw[94] ^ cw[96] ^ cw[98] ^ cw[100] ^ cw[101] ^ cw[104] ^ cw[106] ^ cw[107] ^ cw[110] ^ cw[111] ^ cw[114] ^ cw[115] ^ cw[118] ^ cw[119] ^ cw[121] ^ cw[124] ^ cw[126] ^ cw[128] ^ cw[130] ^ cw[132] ^ cw[134] ^ cw[136] ^ cw[138] ^ cw[140] ^ cw[141] ^ cw[144] ^ cw[145] ^ cw[148] ^ cw[149] ^ cw[152] ^ cw[153] ^ cw[155] ^ cw[158] ^ cw[160] ^ cw[162] ^ cw[164] ^ cw[166] ^ cw[168] ^ cw[170] ^ cw[172] ^ cw[174] ^ cw[176] ^ cw[178] ^ cw[179] ^ cw[182] ^ cw[186] ^ cw[189] ^ cw[192] ^ cw[193] ^ cw[196] ^ cw[199] ^ cw[201] ^ cw[204] ^ cw[206] ^ cw[209] ^ cw[211] ^ cw[213] ^ cw[215] ^ cw[218] ^ cw[220] ^ cw[223] ^ cw[227] ^ cw[228] ^ cw[230] ^ cw[232] ^ cw[235] ^ cw[237] ^ cw[242] ^ cw[245] ^ cw[247] ^ cw[249] ^ cw[251] ^ cw[254] ^ cw[257] ^ cw[259] ^ cw[261] ^ cw[263] ^ cw[267] ^ cw[270] ^ cw[274] ^ cw[277] ^ cw[279] ^ cw[281] ^ cw[283] ^ cw[286] ^ cw[289] ^ cw[290] ^ cw[292] ^ cw[295] ^ cw[296] ^ cw[299] ^ cw[302] ^ cw[305] ^ cw[307] ^ cw[309] ^ cw[310] ^ cw[313] ^ cw[315] ^ cw[316] ^ cw[319] ^ cw[321] ^ cw[323] ^ cw[325] ^ cw[327] ^ cw[329] ^ cw[330] ^ cw[333] ^ cw[335] ^ cw[336] ^ cw[339] ^ cw[341] ^ cw[343] ^ cw[345] ^ cw[347] ^ cw[349] ^ cw[350] ^ cw[353] ^ cw[354] ^ cw[356] ^ cw[358] ^ cw[360] ^ cw[362] ^ cw[364] ^ cw[367] ^ cw[368] ^ cw[371] ^ cw[373] ^ cw[375] ^ cw[377] ^ cw[379] ^ cw[381] ^ cw[383] ^ cw[385] ^ cw[387] ^ cw[389] ^ cw[391] ^ cw[393] ^ cw[394] ^ cw[396] ^ cw[399] ^ cw[401] ^ cw[403] ^ cw[405] ^ cw[407] ^ cw[409] ^ cw[411] ^ cw[413] ^ cw[414] ^ cw[416] ^ cw[419] ^ cw[420] ^ cw[423] ^ cw[424] ^ cw[426] ^ cw[428] ^ cw[430] ^ cw[433] ^ cw[434] ^ cw[437] ^ cw[439] ^ cw[441] ^ cw[443] ^ cw[445] ^ cw[447] ^ cw[449] ^ cw[451] ^ cw[453] ^ cw[455] ^ cw[456] ^ cw[459] ^ cw[460] ^ cw[463] ^ cw[464] ^ cw[466] ^ cw[468] ^ cw[470] ^ cw[473] ^ cw[474] ^ cw[477] ^ cw[478] ^ cw[481] ^ cw[483] ^ cw[485] ^ cw[487] ^ cw[489] ^ cw[491] ^ cw[493] ^ cw[495] ^ cw[496] ^ cw[498] ^ cw[500] ^ cw[502] ^ cw[504] ^ cw[506] ^ cw[508] ^ cw[510] ^ cw[512] ^ cw[515] ^ cw[516] ^ cw[519] ^ cw[521] ^ cw[523] ^ cw[525] ^ cw[527] ^ cw[529] ^ cw[531] ^ cw[533] ^ cw[534] ^ cw[536] ^ cw[538] ^ cw[541] ^ cw[542] ^ cw[545] ^ cw[547] ^ cw[549] ^ cw[551] ^ cw[553] ^ cw[555] ^ cw[557] ^ cw[558] ^ cw[559] ^ cw[561] ^ cw[564] ^ cw[565] ^ cw[568] ^ cw[569] ^ cw[572] ^ cw[573] ^ cw[576] ^ cw[578] ^ cw[579] ^ cw[581] ^ cw[584] ^ cw[586] ^ cw[588] ^ cw[590] ^ cw[592] ^ cw[594] ^ cw[596] ^ cw[598] ^ cw[599] ^ cw[602] ^ cw[603] ^ cw[606] ^ cw[607] ^ cw[610] ^ cw[611] ^ cw[614] ^ cw[616] ^ cw[617] ^ cw[620] ^ cw[621] ^ cw[624] ^ cw[626] ^ cw[628] ^ cw[629] ^ cw[632] ^ cw[633] ^ cw[636] ^ cw[638] ^ cw[639] ^ cw[642] ^ cw[644] ^ cw[646] ^ cw[648] ^ cw[650] ^ cw[652] ^ cw[654] ^ cw[656] ^ cw[657] ^ cw[659] ^ cw[662] ^ cw[663] ^ cw[665] ^ cw[667] ^ cw[669] ^ cw[671] ^ cw[673] ^ cw[676] ^ cw[677] ^ cw[680] ^ cw[681] ^ cw[684] ^ cw[685] ^ cw[688] ^ cw[690] ^ cw[692] ^ cw[694] ^ cw[696] ^ cw[698] ^ cw[699] ^ cw[701] ^ cw[703] ^ cw[706] ^ cw[707] ^ cw[709] ^ cw[711] ^ cw[713] ^ cw[716] ^ cw[717] ^ cw[720] ^ cw[721] ^ cw[724] ^ cw[726] ^ cw[728] ^ cw[730] ^ cw[732] ^ cw[734] ^ cw[736] ^ cw[738] ^ cw[739] ^ cw[742] ^ cw[743] ^ cw[746] ^ cw[747] ^ cw[749] ^ cw[751] ^ cw[753] ^ cw[755] ^ cw[757] ^ cw[759] ^ cw[761] ^ cw[764] ^ cw[765] ^ cw[768] ^ cw[769] ^ cw[772] ^ cw[774] ^ cw[776] ^ cw[778] ^ cw[779] ^ cw[782] ^ cw[783] ^ cw[786] ^ cw[788] ^ cw[789] ^ cw[792] ^ cw[793] ^ cw[796] ^ cw[797] ^ cw[800] ^ cw[801] ^ cw[804] ^ cw[805] ^ cw[808] ^ cw[809] ^ cw[811] ^ cw[813] ^ cw[816] ^ cw[817] ^ cw[819] ^ cw[820] ^ cw[823] ^ cw[824] ^ cw[826] ^ cw[828] ^ cw[830] ^ cw[831] ^ cw[833] ^ cw[835] ^ cw[836] ^ cw[839] ^ cw[841] ^ cw[842] ^ cw[845] ^ cw[847] ^ cw[848] ^ cw[849] ^ cw[851] ^ cw[853] ^ cw[855] ^ cw[856] ^ cw[859] ^ cw[860] ^ cw[861] ^ cw[864] ^ cw[865] ^ cw[866] ^ cw[869] ^ cw[871] ^ cw[872] ^ cw[875] ^ cw[876] ^ cw[878] ^ cw[880] ^ cw[881] ^ cw[883] ^ cw[884] ^ cw[886] ^ cw[888] ^ cw[890] ^ cw[891] ^ cw[893] ^ cw[894] ^ cw[895] ^ cw[897] ^ cw[900] ^ cw[902] ^ cw[904] ^ cw[905] ^ cw[906] ^ cw[908] ^ cw[910] ^ cw[911] ^ cw[914] ^ cw[915] ^ cw[918] ^ cw[920] ^ cw[921] ^ cw[923] ^ cw[925] ^ cw[926] ^ cw[928] ^ cw[929] ^ cw[931] ^ cw[933] ^ cw[935] ^ cw[937] ^ cw[939] ^ cw[941] ^ cw[943] ^ cw[945] ^ cw[947] ^ cw[948] ^ cw[950] ^ cw[952] ^ cw[953] ^ cw[955] ^ cw[956] ^ cw[958] ^ cw[959] ^ cw[961] ^ cw[962] ^ cw[964] ^ cw[965] ^ cw[969] ^ cw[970] ^ cw[971] ^ cw[973] ^ cw[975] ^ cw[976] ^ cw[978] ^ cw[979] ^ cw[980] ^ cw[981] ^ cw[985] ^ cw[986] ^ cw[987] ^ cw[989] ^ cw[991] ^ cw[993] ^ cw[995] ^ cw[997] ^ cw[998] ^ cw[1000] ^ cw[1001] ^ cw[1002] ^ cw[1003] ^ cw[1004] ^ cw[1006] ^ cw[1007] ^ cw[1008] ^ cw[1009] ^ cw[1011] ^ cw[1017];
    assign syndrome[5] = cw[0] ^ cw[2] ^ cw[4] ^ cw[6] ^ cw[8] ^ cw[10] ^ cw[11] ^ cw[13] ^ cw[16] ^ cw[18] ^ cw[20] ^ cw[22] ^ cw[24] ^ cw[26] ^ cw[28] ^ cw[30] ^ cw[32] ^ cw[34] ^ cw[36] ^ cw[38] ^ cw[39] ^ cw[42] ^ cw[44] ^ cw[45] ^ cw[48] ^ cw[50] ^ cw[52] ^ cw[54] ^ cw[56] ^ cw[58] ^ cw[60] ^ cw[62] ^ cw[63] ^ cw[66] ^ cw[68] ^ cw[70] ^ cw[72] ^ cw[73] ^ cw[76] ^ cw[78] ^ cw[80] ^ cw[82] ^ cw[84] ^ cw[86] ^ cw[87] ^ cw[90] ^ cw[91] ^ cw[94] ^ cw[95] ^ cw[97] ^ cw[99] ^ cw[102] ^ cw[103] ^ cw[106] ^ cw[108] ^ cw[110] ^ cw[112] ^ cw[114] ^ cw[116] ^ cw[118] ^ cw[120] ^ cw[121] ^ cw[124] ^ cw[125] ^ cw[128] ^ cw[129] ^ cw[132] ^ cw[133] ^ cw[136] ^ cw[137] ^ cw[140] ^ cw[142] ^ cw[144] ^ cw[146] ^ cw[148] ^ cw[150] ^ cw[151] ^ cw[154] ^ cw[156] ^ cw[158] ^ cw[160] ^ cw[162] ^ cw[164] ^ cw[166] ^ cw[168] ^ cw[170] ^ cw[172] ^ cw[174] ^ cw[175] ^ cw[178] ^ cw[180] ^ cw[182] ^ cw[185] ^ cw[188] ^ cw[191] ^ cw[193] ^ cw[196] ^ cw[198] ^ cw[200] ^ cw[203] ^ cw[206] ^ cw[207] ^ cw[210] ^ cw[213] ^ cw[214] ^ cw[217] ^ cw[222] ^ cw[225] ^ cw[226] ^ cw[229] ^ cw[232] ^ cw[234] ^ cw[236] ^ cw[238] ^ cw[242] ^ cw[245] ^ cw[246] ^ cw[249] ^ cw[252] ^ cw[255] ^ cw[258] ^ cw[259] ^ cw[261] ^ cw[264] ^ cw[267] ^ cw[270] ^ cw[273] ^ cw[276] ^ cw[278] ^ cw[280] ^ cw[284] ^ cw[287] ^ cw[288] ^ cw[289] ^ cw[294] ^ cw[295] ^ cw[298] ^ cw[300] ^ cw[302] ^ cw[304] ^ cw[307] ^ cw[309] ^ cw[311] ^ cw[312] ^ cw[315] ^ cw[317] ^ cw[319] ^ cw[321] ^ cw[323] ^ cw[325] ^ cw[327] ^ cw[329] ^ cw[330] ^ cw[333] ^ cw[334] ^ cw[336] ^ cw[338] ^ cw[340] ^ cw[342] ^ cw[344] ^ cw[346] ^ cw[348] ^ cw[351] ^ cw[352] ^ cw[355] ^ cw[357] ^ cw[359] ^ cw[361] ^ cw[363] ^ cw[365] ^ cw[367] ^ cw[369] ^ cw[371] ^ cw[373] ^ cw[375] ^ cw[377] ^ cw[379] ^ cw[381] ^ cw[383] ^ cw[385] ^ cw[387] ^ cw[389] ^ cw[390] ^ cw[393] ^ cw[395] ^ cw[396] ^ cw[399] ^ cw[400] ^ cw[403] ^ cw[404] ^ cw[407] ^ cw[408] ^ cw[411] ^ cw[412] ^ cw[414] ^ cw[417] ^ cw[418] ^ cw[421] ^ cw[422] ^ cw[425] ^ cw[427] ^ cw[429] ^ cw[431] ^ cw[433] ^ cw[435] ^ cw[437] ^ cw[439] ^ cw[441] ^ cw[443] ^ cw[445] ^ cw[447] ^ cw[449] ^ cw[451] ^ cw[453] ^ cw[455] ^ cw[456] ^ cw[458] ^ cw[460] ^ cw[462] ^ cw[464] ^ cw[467] ^ cw[468] ^ cw[471] ^ cw[472] ^ cw[475] ^ cw[476] ^ cw[479] ^ cw[480] ^ cw[483] ^ cw[484] ^ cw[487] ^ cw[488] ^ cw[491] ^ cw[492] ^ cw[495] ^ cw[497] ^ cw[498] ^ cw[501] ^ cw[502] ^ cw[505] ^ cw[506] ^ cw[509] ^ cw[510] ^ cw[513] ^ cw[514] ^ cw[517] ^ cw[518] ^ cw[521] ^ cw[522] ^ cw[525] ^ cw[526] ^ cw[529] ^ cw[530] ^ cw[533] ^ cw[535] ^ cw[536] ^ cw[539] ^ cw[540] ^ cw[543] ^ cw[544] ^ cw[547] ^ cw[548] ^ cw[551] ^ cw[552] ^ cw[555] ^ cw[556] ^ cw[558] ^ cw[560] ^ cw[562] ^ cw[564] ^ cw[566] ^ cw[568] ^ cw[569] ^ cw[572] ^ cw[574] ^ cw[576] ^ cw[577] ^ cw[579] ^ cw[582] ^ cw[583] ^ cw[586] ^ cw[587] ^ cw[590] ^ cw[591] ^ cw[594] ^ cw[595] ^ cw[598] ^ cw[600] ^ cw[602] ^ cw[604] ^ cw[606] ^ cw[608] ^ cw[609] ^ cw[612] ^ cw[613] ^ cw[616] ^ cw[617] ^ cw[620] ^ cw[621] ^ cw[624] ^ cw[625] ^ cw[628] ^ cw[629] ^ cw[632] ^ cw[633] ^ cw[636] ^ cw[637] ^ cw[639] ^ cw[641] ^ cw[643] ^ cw[645] ^ cw[647] ^ cw[649] ^ cw[651] ^ cw[653] ^ cw[655] ^ cw[658] ^ cw[660] ^ cw[661] ^ cw[664] ^ cw[666] ^ cw[668] ^ cw[670] ^ cw[672] ^ cw[674] ^ cw[676] ^ cw[678] ^ cw[680] ^ cw[682] ^ cw[684] ^ cw[686] ^ cw[688] ^ cw[690] ^ cw[692] ^ cw[694] ^ cw[696] ^ cw[698] ^ cw[699] ^ cw[702] ^ cw[703] ^ cw[706] ^ cw[707] ^ cw[709] ^ cw[711] ^ cw[713] ^ cw[715] ^ cw[717] ^ cw[719] ^ cw[721] ^ cw[723] ^ cw[725] ^ cw[727] ^ cw[729] ^ cw[731] ^ cw[733] ^ cw[735] ^ cw[737] ^ cw[740] ^ cw[741] ^ cw[744] ^ cw[745] ^ cw[748] ^ cw[750] ^ cw[752] ^ cw[754] ^ cw[756] ^ cw[758] ^ cw[760] ^ cw[762] ^ cw[764] ^ cw[766] ^ cw[768] ^ cw[770] ^ cw[772] ^ cw[774] ^ cw[776] ^ cw[778] ^ cw[780] ^ cw[782] ^ cw[784] ^ cw[786] ^ cw[788] ^ cw[789] ^ cw[792] ^ cw[793] ^ cw[796] ^ cw[797] ^ cw[800] ^ cw[801] ^ cw[804] ^ cw[805] ^ cw[808] ^ cw[809] ^ cw[811] ^ cw[812] ^ cw[815] ^ cw[817] ^ cw[818] ^ cw[820] ^ cw[822] ^ cw[824] ^ cw[826] ^ cw[828] ^ cw[829] ^ cw[830] ^ cw[833] ^ cw[834] ^ cw[836] ^ cw[838] ^ cw[840] ^ cw[842] ^ cw[844] ^ cw[845] ^ cw[846] ^ cw[849] ^ cw[851] ^ cw[852] ^ cw[854] ^ cw[857] ^ cw[858] ^ cw[860] ^ cw[862] ^ cw[863] ^ cw[865] ^ cw[867] ^ cw[868] ^ cw[870] ^ cw[873] ^ cw[874] ^ cw[876] ^ cw[878] ^ cw[879] ^ cw[880] ^ cw[882] ^ cw[884] ^ cw[886] ^ cw[887] ^ cw[889] ^ cw[891] ^ cw[893] ^ cw[895] ^ cw[896] ^ cw[898] ^ cw[900] ^ cw[901] ^ cw[904] ^ cw[905] ^ cw[907] ^ cw[909] ^ cw[911] ^ cw[913] ^ cw[914] ^ cw[916] ^ cw[918] ^ cw[920] ^ cw[922] ^ cw[923] ^ cw[924] ^ cw[925] ^ cw[928] ^ cw[930] ^ cw[931] ^ cw[933] ^ cw[935] ^ cw[937] ^ cw[938] ^ cw[940] ^ cw[942] ^ cw[944] ^ cw[946] ^ cw[949] ^ cw[950] ^ cw[951] ^ cw[953] ^ cw[956] ^ cw[957] ^ cw[959] ^ cw[961] ^ cw[963] ^ cw[964] ^ cw[966] ^ cw[967] ^ cw[969] ^ cw[970] ^ cw[971] ^ cw[972] ^ cw[975] ^ cw[976] ^ cw[977] ^ cw[979] ^ cw[981] ^ cw[983] ^ cw[984] ^ cw[986] ^ cw[988] ^ cw[990] ^ cw[992] ^ cw[993] ^ cw[995] ^ cw[996] ^ cw[998] ^ cw[999] ^ cw[1001] ^ cw[1002] ^ cw[1003] ^ cw[1005] ^ cw[1006] ^ cw[1008] ^ cw[1010] ^ cw[1011] ^ cw[1012] ^ cw[1018];
    assign syndrome[4] = cw[0] ^ cw[2] ^ cw[4] ^ cw[6] ^ cw[7] ^ cw[9] ^ cw[12] ^ cw[14] ^ cw[16] ^ cw[18] ^ cw[20] ^ cw[22] ^ cw[24] ^ cw[26] ^ cw[28] ^ cw[30] ^ cw[32] ^ cw[34] ^ cw[35] ^ cw[38] ^ cw[40] ^ cw[41] ^ cw[44] ^ cw[46] ^ cw[48] ^ cw[50] ^ cw[52] ^ cw[54] ^ cw[56] ^ cw[58] ^ cw[60] ^ cw[62] ^ cw[63] ^ cw[66] ^ cw[67] ^ cw[69] ^ cw[71] ^ cw[74] ^ cw[75] ^ cw[78] ^ cw[79] ^ cw[82] ^ cw[83] ^ cw[86] ^ cw[88] ^ cw[90] ^ cw[92] ^ cw[94] ^ cw[96] ^ cw[97] ^ cw[100] ^ cw[101] ^ cw[104] ^ cw[105] ^ cw[108] ^ cw[109] ^ cw[112] ^ cw[113] ^ cw[116] ^ cw[117] ^ cw[120] ^ cw[122] ^ cw[124] ^ cw[126] ^ cw[128] ^ cw[130] ^ cw[132] ^ cw[134] ^ cw[136] ^ cw[138] ^ cw[140] ^ cw[142] ^ cw[144] ^ cw[146] ^ cw[147] ^ cw[150] ^ cw[152] ^ cw[154] ^ cw[156] ^ cw[158] ^ cw[160] ^ cw[162] ^ cw[164] ^ cw[166] ^ cw[168] ^ cw[170] ^ cw[172] ^ cw[174] ^ cw[175] ^ cw[178] ^ cw[179] ^ cw[181] ^ cw[184] ^ cw[187] ^ cw[190] ^ cw[194] ^ cw[196] ^ cw[198] ^ cw[201] ^ cw[202] ^ cw[205] ^ cw[208] ^ cw[210] ^ cw[212] ^ cw[216] ^ cw[219] ^ cw[222] ^ cw[225] ^ cw[226] ^ cw[229] ^ cw[232] ^ cw[234] ^ cw[236] ^ cw[238] ^ cw[242] ^ cw[245] ^ cw[246] ^ cw[249] ^ cw[251] ^ cw[254] ^ cw[257] ^ cw[258] ^ cw[260] ^ cw[263] ^ cw[266] ^ cw[269] ^ cw[272] ^ cw[275] ^ cw[277] ^ cw[279] ^ cw[282] ^ cw[285] ^ cw[287] ^ cw[291] ^ cw[293] ^ cw[295] ^ cw[298] ^ cw[300] ^ cw[302] ^ cw[304] ^ cw[307] ^ cw[309] ^ cw[310] ^ cw[312] ^ cw[314] ^ cw[316] ^ cw[318] ^ cw[320] ^ cw[322] ^ cw[324] ^ cw[326] ^ cw[328] ^ cw[331] ^ cw[332] ^ cw[335] ^ cw[337] ^ cw[339] ^ cw[341] ^ cw[343] ^ cw[345] ^ cw[347] ^ cw[349] ^ cw[351] ^ cw[353] ^ cw[355] ^ cw[357] ^ cw[359] ^ cw[361] ^ cw[363] ^ cw[365] ^ cw[367] ^ cw[369] ^ cw[371] ^ cw[373] ^ cw[375] ^ cw[377] ^ cw[379] ^ cw[381] ^ cw[383] ^ cw[385] ^ cw[387] ^ cw[389] ^ cw[390] ^ cw[393] ^ cw[394] ^ cw[396] ^ cw[398] ^ cw[400] ^ cw[402] ^ cw[404] ^ cw[406] ^ cw[408] ^ cw[410] ^ cw[412] ^ cw[415] ^ cw[416] ^ cw[419] ^ cw[420] ^ cw[423] ^ cw[424] ^ cw[427] ^ cw[428] ^ cw[431] ^ cw[432] ^ cw[435] ^ cw[436] ^ cw[439] ^ cw[440] ^ cw[443] ^ cw[444] ^ cw[447] ^ cw[448] ^ cw[451] ^ cw[452] ^ cw[455] ^ cw[457] ^ cw[458] ^ cw[461] ^ cw[462] ^ cw[465] ^ cw[466] ^ cw[469] ^ cw[470] ^ cw[473] ^ cw[474] ^ cw[477] ^ cw[478] ^ cw[481] ^ cw[482] ^ cw[485] ^ cw[486] ^ cw[489] ^ cw[490] ^ cw[493] ^ cw[494] ^ cw[497] ^ cw[499] ^ cw[501] ^ cw[503] ^ cw[505] ^ cw[507] ^ cw[509] ^ cw[511] ^ cw[513] ^ cw[515] ^ cw[517] ^ cw[519] ^ cw[521] ^ cw[523] ^ cw[525] ^ cw[527] ^ cw[529] ^ cw[531] ^ cw[533] ^ cw[535] ^ cw[536] ^ cw[539] ^ cw[540] ^ cw[543] ^ cw[544] ^ cw[547] ^ cw[548] ^ cw[551] ^ cw[552] ^ cw[555] ^ cw[556] ^ cw[558] ^ cw[559] ^ cw[561] ^ cw[563] ^ cw[565] ^ cw[567] ^ cw[569] ^ cw[571] ^ cw[573] ^ cw[575] ^ cw[577] ^ cw[580] ^ cw[581] ^ cw[584] ^ cw[585] ^ cw[588] ^ cw[589] ^ cw[592] ^ cw[593] ^ cw[596] ^ cw[597] ^ cw[600] ^ cw[601] ^ cw[604] ^ cw[605] ^ cw[608] ^ cw[609] ^ cw[612] ^ cw[613] ^ cw[616] ^ cw[618] ^ cw[620] ^ cw[622] ^ cw[624] ^ cw[625] ^ cw[628] ^ cw[630] ^ cw[632] ^ cw[634] ^ cw[636] ^ cw[638] ^ cw[639] ^ cw[642] ^ cw[643] ^ cw[646] ^ cw[647] ^ cw[650] ^ cw[651] ^ cw[654] ^ cw[655] ^ cw[657] ^ cw[659] ^ cw[662] ^ cw[663] ^ cw[666] ^ cw[667] ^ cw[670] ^ cw[671] ^ cw[674] ^ cw[675] ^ cw[678] ^ cw[679] ^ cw[682] ^ cw[683] ^ cw[686] ^ cw[687] ^ cw[690] ^ cw[691] ^ cw[694] ^ cw[695] ^ cw[698] ^ cw[700] ^ cw[701] ^ cw[704] ^ cw[706] ^ cw[708] ^ cw[709] ^ cw[712] ^ cw[713] ^ cw[716] ^ cw[717] ^ cw[720] ^ cw[721] ^ cw[724] ^ cw[725] ^ cw[728] ^ cw[729] ^ cw[732] ^ cw[733] ^ cw[736] ^ cw[737] ^ cw[740] ^ cw[741] ^ cw[744] ^ cw[745] ^ cw[748] ^ cw[749] ^ cw[752] ^ cw[753] ^ cw[756] ^ cw[757] ^ cw[760] ^ cw[761] ^ cw[764] ^ cw[765] ^ cw[768] ^ cw[769] ^ cw[772] ^ cw[773] ^ cw[776] ^ cw[777] ^ cw[779] ^ cw[781] ^ cw[783] ^ cw[785] ^ cw[787] ^ cw[790] ^ cw[791] ^ cw[794] ^ cw[795] ^ cw[798] ^ cw[799] ^ cw[802] ^ cw[803] ^ cw[806] ^ cw[807] ^ cw[810] ^ cw[812] ^ cw[814] ^ cw[816] ^ cw[817] ^ cw[819] ^ cw[821] ^ cw[823] ^ cw[825] ^ cw[826] ^ cw[828] ^ cw[830] ^ cw[832] ^ cw[833] ^ cw[835] ^ cw[837] ^ cw[839] ^ cw[840] ^ cw[842] ^ cw[845] ^ cw[847] ^ cw[848] ^ cw[849] ^ cw[851] ^ cw[853] ^ cw[855] ^ cw[857] ^ cw[858] ^ cw[860] ^ cw[862] ^ cw[863] ^ cw[864] ^ cw[867] ^ cw[868] ^ cw[870] ^ cw[873] ^ cw[874] ^ cw[876] ^ cw[878] ^ cw[879] ^ cw[881] ^ cw[882] ^ cw[884] ^ cw[886] ^ cw[887] ^ cw[889] ^ cw[890] ^ cw[893] ^ cw[894] ^ cw[897] ^ cw[898] ^ cw[900] ^ cw[901] ^ cw[903] ^ cw[905] ^ cw[906] ^ cw[908] ^ cw[910] ^ cw[912] ^ cw[913] ^ cw[915] ^ cw[917] ^ cw[919] ^ cw[921] ^ cw[924] ^ cw[926] ^ cw[927] ^ cw[929] ^ cw[930] ^ cw[932] ^ cw[934] ^ cw[936] ^ cw[937] ^ cw[939] ^ cw[941] ^ cw[943] ^ cw[945] ^ cw[946] ^ cw[948] ^ cw[950] ^ cw[951] ^ cw[954] ^ cw[956] ^ cw[957] ^ cw[959] ^ cw[961] ^ cw[962] ^ cw[964] ^ cw[965] ^ cw[967] ^ cw[968] ^ cw[969] ^ cw[972] ^ cw[973] ^ cw[974] ^ cw[975] ^ cw[978] ^ cw[980] ^ cw[981] ^ cw[983] ^ cw[984] ^ cw[985] ^ cw[986] ^ cw[987] ^ cw[988] ^ cw[990] ^ cw[991] ^ cw[992] ^ cw[993] ^ cw[994] ^ cw[996] ^ cw[998] ^ cw[1000] ^ cw[1001] ^ cw[1005] ^ cw[1007] ^ cw[1009] ^ cw[1010] ^ cw[1011] ^ cw[1019];
    assign syndrome[3] = cw[0] ^ cw[2] ^ cw[3] ^ cw[5] ^ cw[8] ^ cw[10] ^ cw[12] ^ cw[14] ^ cw[16] ^ cw[18] ^ cw[20] ^ cw[22] ^ cw[24] ^ cw[26] ^ cw[28] ^ cw[30] ^ cw[32] ^ cw[34] ^ cw[35] ^ cw[37] ^ cw[39] ^ cw[42] ^ cw[43] ^ cw[46] ^ cw[47] ^ cw[50] ^ cw[51] ^ cw[54] ^ cw[55] ^ cw[58] ^ cw[59] ^ cw[62] ^ cw[64] ^ cw[66] ^ cw[68] ^ cw[69] ^ cw[72] ^ cw[73] ^ cw[76] ^ cw[77] ^ cw[80] ^ cw[81] ^ cw[84] ^ cw[85] ^ cw[88] ^ cw[89] ^ cw[92] ^ cw[93] ^ cw[96] ^ cw[98] ^ cw[100] ^ cw[102] ^ cw[104] ^ cw[106] ^ cw[108] ^ cw[110] ^ cw[112] ^ cw[114] ^ cw[116] ^ cw[118] ^ cw[120] ^ cw[122] ^ cw[124] ^ cw[126] ^ cw[128] ^ cw[130] ^ cw[132] ^ cw[134] ^ cw[136] ^ cw[138] ^ cw[140] ^ cw[142] ^ cw[144] ^ cw[146] ^ cw[147] ^ cw[150] ^ cw[151] ^ cw[154] ^ cw[155] ^ cw[158] ^ cw[159] ^ cw[162] ^ cw[163] ^ cw[166] ^ cw[167] ^ cw[170] ^ cw[171] ^ cw[174] ^ cw[176] ^ cw[178] ^ cw[180] ^ cw[182] ^ cw[185] ^ cw[188] ^ cw[191] ^ cw[194] ^ cw[195] ^ cw[198] ^ cw[201] ^ cw[203] ^ cw[205] ^ cw[208] ^ cw[209] ^ cw[212] ^ cw[215] ^ cw[218] ^ cw[221] ^ cw[224] ^ cw[225] ^ cw[228] ^ cw[231] ^ cw[233] ^ cw[235] ^ cw[239] ^ cw[241] ^ cw[244] ^ cw[245] ^ cw[247] ^ cw[252] ^ cw[255] ^ cw[258] ^ cw[260] ^ cw[262] ^ cw[265] ^ cw[268] ^ cw[271] ^ cw[274] ^ cw[277] ^ cw[279] ^ cw[281] ^ cw[284] ^ cw[287] ^ cw[289] ^ cw[291] ^ cw[293] ^ cw[295] ^ cw[297] ^ cw[300] ^ cw[302] ^ cw[305] ^ cw[307] ^ cw[309] ^ cw[311] ^ cw[312] ^ cw[315] ^ cw[316] ^ cw[319] ^ cw[320] ^ cw[323] ^ cw[324] ^ cw[327] ^ cw[328] ^ cw[331] ^ cw[332] ^ cw[335] ^ cw[336] ^ cw[339] ^ cw[340] ^ cw[343] ^ cw[344] ^ cw[347] ^ cw[348] ^ cw[351] ^ cw[352] ^ cw[355] ^ cw[356] ^ cw[359] ^ cw[360] ^ cw[363] ^ cw[364] ^ cw[367] ^ cw[368] ^ cw[371] ^ cw[372] ^ cw[375] ^ cw[376] ^ cw[379] ^ cw[380] ^ cw[383] ^ cw[384] ^ cw[387] ^ cw[388] ^ cw[390] ^ cw[392] ^ cw[394] ^ cw[397] ^ cw[398] ^ cw[401] ^ cw[402] ^ cw[405] ^ cw[406] ^ cw[409] ^ cw[410] ^ cw[413] ^ cw[414] ^ cw[417] ^ cw[418] ^ cw[421] ^ cw[422] ^ cw[425] ^ cw[426] ^ cw[429] ^ cw[430] ^ cw[433] ^ cw[434] ^ cw[437] ^ cw[438] ^ cw[441] ^ cw[442] ^ cw[445] ^ cw[446] ^ cw[449] ^ cw[450] ^ cw[453] ^ cw[454] ^ cw[457] ^ cw[459] ^ cw[461] ^ cw[463] ^ cw[465] ^ cw[467] ^ cw[469] ^ cw[471] ^ cw[473] ^ cw[475] ^ cw[477] ^ cw[479] ^ cw[481] ^ cw[483] ^ cw[485] ^ cw[487] ^ cw[489] ^ cw[491] ^ cw[493] ^ cw[495] ^ cw[497] ^ cw[499] ^ cw[501] ^ cw[503] ^ cw[505] ^ cw[507] ^ cw[509] ^ cw[511] ^ cw[513] ^ cw[515] ^ cw[517] ^ cw[519] ^ cw[521] ^ cw[523] ^ cw[525] ^ cw[527] ^ cw[529] ^ cw[531] ^ cw[533] ^ cw[535] ^ cw[536] ^ cw[539] ^ cw[540] ^ cw[543] ^ cw[544] ^ cw[547] ^ cw[548] ^ cw[551] ^ cw[552] ^ cw[555] ^ cw[556] ^ cw[557] ^ cw[559] ^ cw[561] ^ cw[563] ^ cw[565] ^ cw[567] ^ cw[569] ^ cw[571] ^ cw[573] ^ cw[575] ^ cw[577] ^ cw[579] ^ cw[581] ^ cw[583] ^ cw[585] ^ cw[587] ^ cw[589] ^ cw[591] ^ cw[593] ^ cw[595] ^ cw[597] ^ cw[599] ^ cw[601] ^ cw[603] ^ cw[605] ^ cw[607] ^ cw[609] ^ cw[611] ^ cw[613] ^ cw[615] ^ cw[617] ^ cw[619] ^ cw[621] ^ cw[623] ^ cw[625] ^ cw[627] ^ cw[629] ^ cw[631] ^ cw[633] ^ cw[635] ^ cw[637] ^ cw[640] ^ cw[641] ^ cw[644] ^ cw[645] ^ cw[648] ^ cw[649] ^ cw[652] ^ cw[653] ^ cw[656] ^ cw[657] ^ cw[660] ^ cw[661] ^ cw[664] ^ cw[665] ^ cw[668] ^ cw[669] ^ cw[672] ^ cw[673] ^ cw[676] ^ cw[677] ^ cw[680] ^ cw[681] ^ cw[684] ^ cw[685] ^ cw[688] ^ cw[689] ^ cw[692] ^ cw[693] ^ cw[696] ^ cw[697] ^ cw[700] ^ cw[701] ^ cw[704] ^ cw[705] ^ cw[708] ^ cw[710] ^ cw[712] ^ cw[714] ^ cw[716] ^ cw[718] ^ cw[720] ^ cw[722] ^ cw[724] ^ cw[726] ^ cw[728] ^ cw[730] ^ cw[732] ^ cw[734] ^ cw[736] ^ cw[738] ^ cw[740] ^ cw[742] ^ cw[744] ^ cw[746] ^ cw[748] ^ cw[750] ^ cw[752] ^ cw[754] ^ cw[756] ^ cw[758] ^ cw[760] ^ cw[762] ^ cw[764] ^ cw[766] ^ cw[768] ^ cw[770] ^ cw[772] ^ cw[774] ^ cw[776] ^ cw[778] ^ cw[779] ^ cw[782] ^ cw[783] ^ cw[786] ^ cw[787] ^ cw[790] ^ cw[791] ^ cw[794] ^ cw[795] ^ cw[798] ^ cw[799] ^ cw[802] ^ cw[803] ^ cw[806] ^ cw[807] ^ cw[810] ^ cw[811] ^ cw[813] ^ cw[814] ^ cw[816] ^ cw[819] ^ cw[820] ^ cw[823] ^ cw[824] ^ cw[826] ^ cw[827] ^ cw[830] ^ cw[831] ^ cw[832] ^ cw[834] ^ cw[836] ^ cw[838] ^ cw[840] ^ cw[841] ^ cw[843] ^ cw[844] ^ cw[846] ^ cw[848] ^ cw[850] ^ cw[852] ^ cw[854] ^ cw[856] ^ cw[857] ^ cw[859] ^ cw[861] ^ cw[862] ^ cw[865] ^ cw[866] ^ cw[868] ^ cw[869] ^ cw[871] ^ cw[872] ^ cw[874] ^ cw[876] ^ cw[877] ^ cw[878] ^ cw[881] ^ cw[883] ^ cw[885] ^ cw[886] ^ cw[888] ^ cw[891] ^ cw[892] ^ cw[893] ^ cw[895] ^ cw[898] ^ cw[899] ^ cw[901] ^ cw[904] ^ cw[905] ^ cw[907] ^ cw[909] ^ cw[910] ^ cw[913] ^ cw[914] ^ cw[916] ^ cw[918] ^ cw[920] ^ cw[921] ^ cw[922] ^ cw[924] ^ cw[926] ^ cw[927] ^ cw[930] ^ cw[932] ^ cw[934] ^ cw[936] ^ cw[937] ^ cw[939] ^ cw[941] ^ cw[943] ^ cw[945] ^ cw[946] ^ cw[948] ^ cw[949] ^ cw[951] ^ cw[953] ^ cw[954] ^ cw[956] ^ cw[959] ^ cw[961] ^ cw[962] ^ cw[963] ^ cw[964] ^ cw[965] ^ cw[966] ^ cw[968] ^ cw[971] ^ cw[973] ^ cw[974] ^ cw[976] ^ cw[977] ^ cw[979] ^ cw[982] ^ cw[983] ^ cw[985] ^ cw[986] ^ cw[989] ^ cw[990] ^ cw[992] ^ cw[993] ^ cw[995] ^ cw[996] ^ cw[997] ^ cw[999] ^ cw[1000] ^ cw[1002] ^ cw[1003] ^ cw[1004] ^ cw[1005] ^ cw[1006] ^ cw[1008] ^ cw[1010] ^ cw[1012] ^ cw[1020];
    assign syndrome[2] = cw[0] ^ cw[1] ^ cw[3] ^ cw[6] ^ cw[7] ^ cw[10] ^ cw[11] ^ cw[14] ^ cw[15] ^ cw[18] ^ cw[19] ^ cw[22] ^ cw[23] ^ cw[26] ^ cw[27] ^ cw[30] ^ cw[31] ^ cw[34] ^ cw[36] ^ cw[37] ^ cw[40] ^ cw[41] ^ cw[44] ^ cw[45] ^ cw[48] ^ cw[49] ^ cw[52] ^ cw[53] ^ cw[56] ^ cw[57] ^ cw[60] ^ cw[61] ^ cw[64] ^ cw[65] ^ cw[68] ^ cw[70] ^ cw[72] ^ cw[74] ^ cw[76] ^ cw[78] ^ cw[80] ^ cw[82] ^ cw[84] ^ cw[86] ^ cw[88] ^ cw[90] ^ cw[92] ^ cw[94] ^ cw[96] ^ cw[98] ^ cw[100] ^ cw[102] ^ cw[104] ^ cw[106] ^ cw[108] ^ cw[110] ^ cw[112] ^ cw[114] ^ cw[116] ^ cw[118] ^ cw[120] ^ cw[122] ^ cw[124] ^ cw[126] ^ cw[128] ^ cw[130] ^ cw[132] ^ cw[134] ^ cw[136] ^ cw[138] ^ cw[140] ^ cw[142] ^ cw[144] ^ cw[146] ^ cw[147] ^ cw[150] ^ cw[151] ^ cw[154] ^ cw[155] ^ cw[158] ^ cw[159] ^ cw[162] ^ cw[163] ^ cw[166] ^ cw[167] ^ cw[170] ^ cw[171] ^ cw[174] ^ cw[175] ^ cw[178] ^ cw[179] ^ cw[181] ^ cw[184] ^ cw[187] ^ cw[190] ^ cw[193] ^ cw[195] ^ cw[197] ^ cw[200] ^ cw[202] ^ cw[204] ^ cw[207] ^ cw[209] ^ cw[211] ^ cw[214] ^ cw[217] ^ cw[220] ^ cw[223] ^ cw[225] ^ cw[227] ^ cw[230] ^ cw[232] ^ cw[234] ^ cw[237] ^ cw[240] ^ cw[243] ^ cw[245] ^ cw[248] ^ cw[250] ^ cw[253] ^ cw[256] ^ cw[258] ^ cw[262] ^ cw[265] ^ cw[268] ^ cw[271] ^ cw[274] ^ cw[277] ^ cw[279] ^ cw[281] ^ cw[284] ^ cw[287] ^ cw[289] ^ cw[291] ^ cw[293] ^ cw[295] ^ cw[297] ^ cw[300] ^ cw[302] ^ cw[304] ^ cw[307] ^ cw[309] ^ cw[310] ^ cw[312] ^ cw[314] ^ cw[316] ^ cw[318] ^ cw[320] ^ cw[322] ^ cw[324] ^ cw[326] ^ cw[328] ^ cw[330] ^ cw[332] ^ cw[334] ^ cw[336] ^ cw[338] ^ cw[340] ^ cw[342] ^ cw[344] ^ cw[346] ^ cw[348] ^ cw[350] ^ cw[352] ^ cw[354] ^ cw[356] ^ cw[358] ^ cw[360] ^ cw[362] ^ cw[364] ^ cw[366] ^ cw[368] ^ cw[370] ^ cw[372] ^ cw[374] ^ cw[376] ^ cw[378] ^ cw[380] ^ cw[382] ^ cw[384] ^ cw[386] ^ cw[388] ^ cw[391] ^ cw[392] ^ cw[395] ^ cw[396] ^ cw[399] ^ cw[400] ^ cw[403] ^ cw[404] ^ cw[407] ^ cw[408] ^ cw[411] ^ cw[412] ^ cw[415] ^ cw[416] ^ cw[419] ^ cw[420] ^ cw[423] ^ cw[424] ^ cw[427] ^ cw[428] ^ cw[431] ^ cw[432] ^ cw[435] ^ cw[436] ^ cw[439] ^ cw[440] ^ cw[443] ^ cw[444] ^ cw[447] ^ cw[448] ^ cw[451] ^ cw[452] ^ cw[455] ^ cw[456] ^ cw[459] ^ cw[460] ^ cw[463] ^ cw[464] ^ cw[467] ^ cw[468] ^ cw[471] ^ cw[472] ^ cw[475] ^ cw[476] ^ cw[479] ^ cw[480] ^ cw[483] ^ cw[484] ^ cw[487] ^ cw[488] ^ cw[491] ^ cw[492] ^ cw[495] ^ cw[496] ^ cw[499] ^ cw[500] ^ cw[503] ^ cw[504] ^ cw[507] ^ cw[508] ^ cw[511] ^ cw[512] ^ cw[515] ^ cw[516] ^ cw[519] ^ cw[520] ^ cw[523] ^ cw[524] ^ cw[527] ^ cw[528] ^ cw[531] ^ cw[532] ^ cw[535] ^ cw[537] ^ cw[539] ^ cw[541] ^ cw[543] ^ cw[545] ^ cw[547] ^ cw[549] ^ cw[551] ^ cw[553] ^ cw[555] ^ cw[556] ^ cw[558] ^ cw[559] ^ cw[562] ^ cw[563] ^ cw[566] ^ cw[567] ^ cw[568] ^ cw[571] ^ cw[574] ^ cw[575] ^ cw[576] ^ cw[579] ^ cw[582] ^ cw[583] ^ cw[586] ^ cw[587] ^ cw[590] ^ cw[591] ^ cw[594] ^ cw[595] ^ cw[598] ^ cw[599] ^ cw[602] ^ cw[603] ^ cw[606] ^ cw[607] ^ cw[608] ^ cw[611] ^ cw[612] ^ cw[615] ^ cw[618] ^ cw[619] ^ cw[622] ^ cw[623] ^ cw[624] ^ cw[627] ^ cw[630] ^ cw[631] ^ cw[634] ^ cw[635] ^ cw[638] ^ cw[639] ^ cw[642] ^ cw[643] ^ cw[646] ^ cw[647] ^ cw[650] ^ cw[651] ^ cw[654] ^ cw[655] ^ cw[656] ^ cw[659] ^ cw[662] ^ cw[663] ^ cw[666] ^ cw[667] ^ cw[670] ^ cw[671] ^ cw[674] ^ cw[675] ^ cw[678] ^ cw[679] ^ cw[682] ^ cw[683] ^ cw[686] ^ cw[687] ^ cw[690] ^ cw[691] ^ cw[694] ^ cw[695] ^ cw[698] ^ cw[699] ^ cw[700] ^ cw[703] ^ cw[706] ^ cw[707] ^ cw[710] ^ cw[711] ^ cw[714] ^ cw[715] ^ cw[718] ^ cw[719] ^ cw[722] ^ cw[723] ^ cw[726] ^ cw[727] ^ cw[730] ^ cw[731] ^ cw[734] ^ cw[735] ^ cw[738] ^ cw[739] ^ cw[742] ^ cw[743] ^ cw[746] ^ cw[747] ^ cw[750] ^ cw[751] ^ cw[754] ^ cw[755] ^ cw[758] ^ cw[759] ^ cw[762] ^ cw[763] ^ cw[766] ^ cw[767] ^ cw[770] ^ cw[771] ^ cw[774] ^ cw[775] ^ cw[778] ^ cw[780] ^ cw[782] ^ cw[784] ^ cw[786] ^ cw[788] ^ cw[790] ^ cw[792] ^ cw[794] ^ cw[796] ^ cw[798] ^ cw[800] ^ cw[802] ^ cw[804] ^ cw[806] ^ cw[808] ^ cw[810] ^ cw[812] ^ cw[814] ^ cw[816] ^ cw[818] ^ cw[819] ^ cw[821] ^ cw[823] ^ cw[825] ^ cw[826] ^ cw[827] ^ cw[829] ^ cw[832] ^ cw[833] ^ cw[835] ^ cw[837] ^ cw[839] ^ cw[840] ^ cw[841] ^ cw[843] ^ cw[845] ^ cw[847] ^ cw[850] ^ cw[851] ^ cw[853] ^ cw[855] ^ cw[857] ^ cw[859] ^ cw[860] ^ cw[862] ^ cw[864] ^ cw[865] ^ cw[867] ^ cw[868] ^ cw[869] ^ cw[871] ^ cw[873] ^ cw[874] ^ cw[875] ^ cw[878] ^ cw[880] ^ cw[883] ^ cw[884] ^ cw[886] ^ cw[888] ^ cw[889] ^ cw[891] ^ cw[893] ^ cw[895] ^ cw[896] ^ cw[898] ^ cw[900] ^ cw[901] ^ cw[902] ^ cw[904] ^ cw[907] ^ cw[909] ^ cw[910] ^ cw[911] ^ cw[913] ^ cw[916] ^ cw[918] ^ cw[920] ^ cw[921] ^ cw[922] ^ cw[924] ^ cw[926] ^ cw[929] ^ cw[930] ^ cw[932] ^ cw[934] ^ cw[936] ^ cw[937] ^ cw[939] ^ cw[941] ^ cw[943] ^ cw[945] ^ cw[946] ^ cw[948] ^ cw[949] ^ cw[951] ^ cw[953] ^ cw[954] ^ cw[957] ^ cw[959] ^ cw[961] ^ cw[962] ^ cw[963] ^ cw[965] ^ cw[966] ^ cw[968] ^ cw[969] ^ cw[971] ^ cw[972] ^ cw[974] ^ cw[975] ^ cw[976] ^ cw[977] ^ cw[979] ^ cw[980] ^ cw[981] ^ cw[982] ^ cw[984] ^ cw[985] ^ cw[987] ^ cw[988] ^ cw[989] ^ cw[991] ^ cw[992] ^ cw[994] ^ cw[996] ^ cw[997] ^ cw[999] ^ cw[1003] ^ cw[1004] ^ cw[1006] ^ cw[1007] ^ cw[1009] ^ cw[1012] ^ cw[1021];
    assign syndrome[1] = cw[0] ^ cw[1] ^ cw[3] ^ cw[5] ^ cw[7] ^ cw[9] ^ cw[11] ^ cw[13] ^ cw[15] ^ cw[17] ^ cw[19] ^ cw[21] ^ cw[23] ^ cw[25] ^ cw[27] ^ cw[29] ^ cw[31] ^ cw[33] ^ cw[35] ^ cw[38] ^ cw[39] ^ cw[42] ^ cw[43] ^ cw[46] ^ cw[47] ^ cw[50] ^ cw[51] ^ cw[54] ^ cw[55] ^ cw[58] ^ cw[59] ^ cw[62] ^ cw[63] ^ cw[66] ^ cw[67] ^ cw[70] ^ cw[71] ^ cw[74] ^ cw[75] ^ cw[78] ^ cw[79] ^ cw[82] ^ cw[83] ^ cw[86] ^ cw[87] ^ cw[90] ^ cw[91] ^ cw[94] ^ cw[95] ^ cw[98] ^ cw[99] ^ cw[102] ^ cw[103] ^ cw[106] ^ cw[107] ^ cw[110] ^ cw[111] ^ cw[114] ^ cw[115] ^ cw[118] ^ cw[119] ^ cw[122] ^ cw[123] ^ cw[126] ^ cw[127] ^ cw[130] ^ cw[131] ^ cw[134] ^ cw[135] ^ cw[138] ^ cw[139] ^ cw[142] ^ cw[143] ^ cw[146] ^ cw[148] ^ cw[150] ^ cw[152] ^ cw[154] ^ cw[156] ^ cw[158] ^ cw[160] ^ cw[162] ^ cw[164] ^ cw[166] ^ cw[168] ^ cw[170] ^ cw[172] ^ cw[174] ^ cw[176] ^ cw[178] ^ cw[180] ^ cw[183] ^ cw[186] ^ cw[189] ^ cw[192] ^ cw[195] ^ cw[197] ^ cw[199] ^ cw[202] ^ cw[204] ^ cw[206] ^ cw[209] ^ cw[211] ^ cw[213] ^ cw[216] ^ cw[219] ^ cw[222] ^ cw[225] ^ cw[227] ^ cw[229] ^ cw[232] ^ cw[234] ^ cw[236] ^ cw[239] ^ cw[242] ^ cw[245] ^ cw[247] ^ cw[249] ^ cw[252] ^ cw[255] ^ cw[258] ^ cw[260] ^ cw[262] ^ cw[265] ^ cw[268] ^ cw[271] ^ cw[274] ^ cw[277] ^ cw[279] ^ cw[281] ^ cw[284] ^ cw[287] ^ cw[289] ^ cw[291] ^ cw[293] ^ cw[294] ^ cw[297] ^ cw[298] ^ cw[302] ^ cw[304] ^ cw[305] ^ cw[309] ^ cw[310] ^ cw[312] ^ cw[314] ^ cw[316] ^ cw[318] ^ cw[320] ^ cw[322] ^ cw[324] ^ cw[326] ^ cw[328] ^ cw[330] ^ cw[332] ^ cw[334] ^ cw[336] ^ cw[338] ^ cw[340] ^ cw[342] ^ cw[344] ^ cw[346] ^ cw[348] ^ cw[350] ^ cw[352] ^ cw[354] ^ cw[356] ^ cw[358] ^ cw[360] ^ cw[362] ^ cw[364] ^ cw[366] ^ cw[368] ^ cw[370] ^ cw[372] ^ cw[374] ^ cw[376] ^ cw[378] ^ cw[380] ^ cw[382] ^ cw[384] ^ cw[386] ^ cw[388] ^ cw[390] ^ cw[392] ^ cw[394] ^ cw[396] ^ cw[398] ^ cw[400] ^ cw[402] ^ cw[404] ^ cw[406] ^ cw[408] ^ cw[410] ^ cw[412] ^ cw[414] ^ cw[416] ^ cw[418] ^ cw[420] ^ cw[422] ^ cw[424] ^ cw[426] ^ cw[428] ^ cw[430] ^ cw[432] ^ cw[434] ^ cw[436] ^ cw[438] ^ cw[440] ^ cw[442] ^ cw[444] ^ cw[446] ^ cw[448] ^ cw[450] ^ cw[452] ^ cw[454] ^ cw[456] ^ cw[458] ^ cw[460] ^ cw[462] ^ cw[464] ^ cw[466] ^ cw[468] ^ cw[470] ^ cw[472] ^ cw[474] ^ cw[476] ^ cw[478] ^ cw[480] ^ cw[482] ^ cw[484] ^ cw[486] ^ cw[488] ^ cw[490] ^ cw[492] ^ cw[494] ^ cw[496] ^ cw[498] ^ cw[500] ^ cw[502] ^ cw[504] ^ cw[506] ^ cw[508] ^ cw[510] ^ cw[512] ^ cw[514] ^ cw[516] ^ cw[518] ^ cw[520] ^ cw[522] ^ cw[524] ^ cw[526] ^ cw[528] ^ cw[530] ^ cw[532] ^ cw[534] ^ cw[536] ^ cw[538] ^ cw[540] ^ cw[542] ^ cw[544] ^ cw[546] ^ cw[548] ^ cw[550] ^ cw[552] ^ cw[554] ^ cw[555] ^ cw[558] ^ cw[560] ^ cw[561] ^ cw[564] ^ cw[565] ^ cw[568] ^ cw[570] ^ cw[572] ^ cw[573] ^ cw[576] ^ cw[578] ^ cw[580] ^ cw[581] ^ cw[584] ^ cw[585] ^ cw[588] ^ cw[589] ^ cw[592] ^ cw[593] ^ cw[596] ^ cw[597] ^ cw[600] ^ cw[601] ^ cw[604] ^ cw[605] ^ cw[608] ^ cw[610] ^ cw[612] ^ cw[614] ^ cw[616] ^ cw[617] ^ cw[620] ^ cw[621] ^ cw[624] ^ cw[626] ^ cw[628] ^ cw[629] ^ cw[632] ^ cw[633] ^ cw[636] ^ cw[637] ^ cw[640] ^ cw[641] ^ cw[644] ^ cw[645] ^ cw[648] ^ cw[649] ^ cw[652] ^ cw[653] ^ cw[656] ^ cw[658] ^ cw[660] ^ cw[661] ^ cw[664] ^ cw[665] ^ cw[668] ^ cw[669] ^ cw[672] ^ cw[673] ^ cw[676] ^ cw[677] ^ cw[680] ^ cw[681] ^ cw[684] ^ cw[685] ^ cw[688] ^ cw[689] ^ cw[692] ^ cw[693] ^ cw[696] ^ cw[697] ^ cw[700] ^ cw[702] ^ cw[704] ^ cw[705] ^ cw[708] ^ cw[709] ^ cw[712] ^ cw[713] ^ cw[716] ^ cw[717] ^ cw[720] ^ cw[721] ^ cw[724] ^ cw[725] ^ cw[728] ^ cw[729] ^ cw[732] ^ cw[733] ^ cw[736] ^ cw[737] ^ cw[740] ^ cw[741] ^ cw[744] ^ cw[745] ^ cw[748] ^ cw[749] ^ cw[752] ^ cw[753] ^ cw[756] ^ cw[757] ^ cw[760] ^ cw[761] ^ cw[764] ^ cw[765] ^ cw[768] ^ cw[769] ^ cw[772] ^ cw[773] ^ cw[776] ^ cw[777] ^ cw[780] ^ cw[781] ^ cw[784] ^ cw[785] ^ cw[788] ^ cw[789] ^ cw[792] ^ cw[793] ^ cw[796] ^ cw[797] ^ cw[800] ^ cw[801] ^ cw[804] ^ cw[805] ^ cw[808] ^ cw[809] ^ cw[812] ^ cw[814] ^ cw[815] ^ cw[818] ^ cw[819] ^ cw[821] ^ cw[822] ^ cw[825] ^ cw[827] ^ cw[829] ^ cw[830] ^ cw[832] ^ cw[833] ^ cw[835] ^ cw[837] ^ cw[839] ^ cw[841] ^ cw[843] ^ cw[845] ^ cw[847] ^ cw[848] ^ cw[850] ^ cw[851] ^ cw[853] ^ cw[855] ^ cw[857] ^ cw[859] ^ cw[860] ^ cw[862] ^ cw[864] ^ cw[865] ^ cw[867] ^ cw[869] ^ cw[871] ^ cw[873] ^ cw[875] ^ cw[876] ^ cw[878] ^ cw[880] ^ cw[881] ^ cw[883] ^ cw[884] ^ cw[886] ^ cw[888] ^ cw[889] ^ cw[891] ^ cw[893] ^ cw[895] ^ cw[896] ^ cw[898] ^ cw[900] ^ cw[902] ^ cw[904] ^ cw[905] ^ cw[907] ^ cw[909] ^ cw[911] ^ cw[913] ^ cw[914] ^ cw[916] ^ cw[918] ^ cw[920] ^ cw[922] ^ cw[924] ^ cw[926] ^ cw[927] ^ cw[929] ^ cw[930] ^ cw[932] ^ cw[934] ^ cw[936] ^ cw[937] ^ cw[939] ^ cw[941] ^ cw[943] ^ cw[945] ^ cw[946] ^ cw[948] ^ cw[949] ^ cw[951] ^ cw[953] ^ cw[954] ^ cw[956] ^ cw[957] ^ cw[959] ^ cw[962] ^ cw[963] ^ cw[964] ^ cw[965] ^ cw[966] ^ cw[968] ^ cw[969] ^ cw[971] ^ cw[973] ^ cw[974] ^ cw[976] ^ cw[977] ^ cw[979] ^ cw[980] ^ cw[981] ^ cw[983] ^ cw[984] ^ cw[986] ^ cw[987] ^ cw[988] ^ cw[990] ^ cw[991] ^ cw[993] ^ cw[994] ^ cw[995] ^ cw[999] ^ cw[1000] ^ cw[1002] ^ cw[1004] ^ cw[1005] ^ cw[1008] ^ cw[1010] ^ cw[1012] ^ cw[1022];
    assign syndrome[0] = cw[0] ^ cw[1] ^ cw[2] ^ cw[5] ^ cw[6] ^ cw[9] ^ cw[10] ^ cw[13] ^ cw[14] ^ cw[17] ^ cw[18] ^ cw[21] ^ cw[22] ^ cw[25] ^ cw[26] ^ cw[29] ^ cw[30] ^ cw[33] ^ cw[34] ^ cw[37] ^ cw[38] ^ cw[41] ^ cw[42] ^ cw[45] ^ cw[46] ^ cw[49] ^ cw[50] ^ cw[53] ^ cw[54] ^ cw[57] ^ cw[58] ^ cw[61] ^ cw[62] ^ cw[65] ^ cw[66] ^ cw[69] ^ cw[70] ^ cw[73] ^ cw[74] ^ cw[77] ^ cw[78] ^ cw[81] ^ cw[82] ^ cw[85] ^ cw[86] ^ cw[89] ^ cw[90] ^ cw[93] ^ cw[94] ^ cw[97] ^ cw[98] ^ cw[101] ^ cw[102] ^ cw[105] ^ cw[106] ^ cw[109] ^ cw[110] ^ cw[113] ^ cw[114] ^ cw[117] ^ cw[118] ^ cw[121] ^ cw[122] ^ cw[125] ^ cw[126] ^ cw[129] ^ cw[130] ^ cw[133] ^ cw[134] ^ cw[137] ^ cw[138] ^ cw[141] ^ cw[142] ^ cw[145] ^ cw[146] ^ cw[149] ^ cw[150] ^ cw[153] ^ cw[154] ^ cw[157] ^ cw[158] ^ cw[161] ^ cw[162] ^ cw[165] ^ cw[166] ^ cw[169] ^ cw[170] ^ cw[173] ^ cw[174] ^ cw[177] ^ cw[178] ^ cw[183] ^ cw[186] ^ cw[189] ^ cw[192] ^ cw[195] ^ cw[197] ^ cw[199] ^ cw[202] ^ cw[204] ^ cw[206] ^ cw[209] ^ cw[211] ^ cw[213] ^ cw[216] ^ cw[219] ^ cw[222] ^ cw[225] ^ cw[227] ^ cw[229] ^ cw[232] ^ cw[234] ^ cw[236] ^ cw[239] ^ cw[242] ^ cw[245] ^ cw[247] ^ cw[249] ^ cw[252] ^ cw[255] ^ cw[258] ^ cw[260] ^ cw[262] ^ cw[265] ^ cw[268] ^ cw[271] ^ cw[274] ^ cw[277] ^ cw[279] ^ cw[281] ^ cw[284] ^ cw[287] ^ cw[289] ^ cw[291] ^ cw[293] ^ cw[294] ^ cw[297] ^ cw[298] ^ cw[300] ^ cw[304] ^ cw[305] ^ cw[307] ^ cw[310] ^ cw[311] ^ cw[314] ^ cw[315] ^ cw[318] ^ cw[319] ^ cw[322] ^ cw[323] ^ cw[326] ^ cw[327] ^ cw[330] ^ cw[331] ^ cw[334] ^ cw[335] ^ cw[338] ^ cw[339] ^ cw[342] ^ cw[343] ^ cw[346] ^ cw[347] ^ cw[350] ^ cw[351] ^ cw[354] ^ cw[355] ^ cw[358] ^ cw[359] ^ cw[362] ^ cw[363] ^ cw[366] ^ cw[367] ^ cw[370] ^ cw[371] ^ cw[374] ^ cw[375] ^ cw[378] ^ cw[379] ^ cw[382] ^ cw[383] ^ cw[386] ^ cw[387] ^ cw[390] ^ cw[391] ^ cw[394] ^ cw[395] ^ cw[398] ^ cw[399] ^ cw[402] ^ cw[403] ^ cw[406] ^ cw[407] ^ cw[410] ^ cw[411] ^ cw[414] ^ cw[415] ^ cw[418] ^ cw[419] ^ cw[422] ^ cw[423] ^ cw[426] ^ cw[427] ^ cw[430] ^ cw[431] ^ cw[434] ^ cw[435] ^ cw[438] ^ cw[439] ^ cw[442] ^ cw[443] ^ cw[446] ^ cw[447] ^ cw[450] ^ cw[451] ^ cw[454] ^ cw[455] ^ cw[458] ^ cw[459] ^ cw[462] ^ cw[463] ^ cw[466] ^ cw[467] ^ cw[470] ^ cw[471] ^ cw[474] ^ cw[475] ^ cw[478] ^ cw[479] ^ cw[482] ^ cw[483] ^ cw[486] ^ cw[487] ^ cw[490] ^ cw[491] ^ cw[494] ^ cw[495] ^ cw[498] ^ cw[499] ^ cw[502] ^ cw[503] ^ cw[506] ^ cw[507] ^ cw[510] ^ cw[511] ^ cw[514] ^ cw[515] ^ cw[518] ^ cw[519] ^ cw[522] ^ cw[523] ^ cw[526] ^ cw[527] ^ cw[530] ^ cw[531] ^ cw[534] ^ cw[535] ^ cw[538] ^ cw[539] ^ cw[542] ^ cw[543] ^ cw[546] ^ cw[547] ^ cw[550] ^ cw[551] ^ cw[554] ^ cw[556] ^ cw[557] ^ cw[559] ^ cw[560] ^ cw[563] ^ cw[564] ^ cw[567] ^ cw[569] ^ cw[571] ^ cw[572] ^ cw[575] ^ cw[577] ^ cw[579] ^ cw[580] ^ cw[583] ^ cw[584] ^ cw[587] ^ cw[588] ^ cw[591] ^ cw[592] ^ cw[595] ^ cw[596] ^ cw[599] ^ cw[600] ^ cw[603] ^ cw[604] ^ cw[607] ^ cw[609] ^ cw[611] ^ cw[613] ^ cw[615] ^ cw[616] ^ cw[619] ^ cw[620] ^ cw[623] ^ cw[625] ^ cw[627] ^ cw[628] ^ cw[631] ^ cw[632] ^ cw[635] ^ cw[636] ^ cw[639] ^ cw[640] ^ cw[643] ^ cw[644] ^ cw[647] ^ cw[648] ^ cw[651] ^ cw[652] ^ cw[655] ^ cw[657] ^ cw[659] ^ cw[660] ^ cw[663] ^ cw[664] ^ cw[667] ^ cw[668] ^ cw[671] ^ cw[672] ^ cw[675] ^ cw[676] ^ cw[679] ^ cw[680] ^ cw[683] ^ cw[684] ^ cw[687] ^ cw[688] ^ cw[691] ^ cw[692] ^ cw[695] ^ cw[696] ^ cw[699] ^ cw[701] ^ cw[703] ^ cw[704] ^ cw[707] ^ cw[708] ^ cw[711] ^ cw[712] ^ cw[715] ^ cw[716] ^ cw[719] ^ cw[720] ^ cw[723] ^ cw[724] ^ cw[727] ^ cw[728] ^ cw[731] ^ cw[732] ^ cw[735] ^ cw[736] ^ cw[739] ^ cw[740] ^ cw[743] ^ cw[744] ^ cw[747] ^ cw[748] ^ cw[751] ^ cw[752] ^ cw[755] ^ cw[756] ^ cw[759] ^ cw[760] ^ cw[763] ^ cw[764] ^ cw[767] ^ cw[768] ^ cw[771] ^ cw[772] ^ cw[775] ^ cw[776] ^ cw[779] ^ cw[780] ^ cw[783] ^ cw[784] ^ cw[787] ^ cw[788] ^ cw[791] ^ cw[792] ^ cw[795] ^ cw[796] ^ cw[799] ^ cw[800] ^ cw[803] ^ cw[804] ^ cw[807] ^ cw[808] ^ cw[811] ^ cw[813] ^ cw[814] ^ cw[817] ^ cw[818] ^ cw[820] ^ cw[821] ^ cw[824] ^ cw[825] ^ cw[828] ^ cw[829] ^ cw[831] ^ cw[832] ^ cw[834] ^ cw[836] ^ cw[838] ^ cw[839] ^ cw[842] ^ cw[843] ^ cw[844] ^ cw[846] ^ cw[849] ^ cw[850] ^ cw[852] ^ cw[854] ^ cw[856] ^ cw[858] ^ cw[859] ^ cw[861] ^ cw[863] ^ cw[864] ^ cw[866] ^ cw[867] ^ cw[870] ^ cw[871] ^ cw[872] ^ cw[873] ^ cw[875] ^ cw[877] ^ cw[879] ^ cw[882] ^ cw[883] ^ cw[885] ^ cw[887] ^ cw[888] ^ cw[890] ^ cw[892] ^ cw[894] ^ cw[895] ^ cw[897] ^ cw[899] ^ cw[900] ^ cw[903] ^ cw[904] ^ cw[906] ^ cw[908] ^ cw[909] ^ cw[912] ^ cw[913] ^ cw[915] ^ cw[917] ^ cw[919] ^ cw[920] ^ cw[922] ^ cw[923] ^ cw[925] ^ cw[928] ^ cw[929] ^ cw[931] ^ cw[933] ^ cw[935] ^ cw[936] ^ cw[938] ^ cw[940] ^ cw[942] ^ cw[944] ^ cw[945] ^ cw[947] ^ cw[949] ^ cw[950] ^ cw[952] ^ cw[954] ^ cw[955] ^ cw[957] ^ cw[958] ^ cw[960] ^ cw[961] ^ cw[963] ^ cw[965] ^ cw[966] ^ cw[967] ^ cw[969] ^ cw[970] ^ cw[972] ^ cw[974] ^ cw[975] ^ cw[977] ^ cw[978] ^ cw[980] ^ cw[981] ^ cw[982] ^ cw[984] ^ cw[985] ^ cw[987] ^ cw[988] ^ cw[989] ^ cw[991] ^ cw[992] ^ cw[994] ^ cw[996] ^ cw[997] ^ cw[998] ^ cw[1001] ^ cw[1003] ^ cw[1006] ^ cw[1007] ^ cw[1009] ^ cw[1011] ^ cw[1023];
    assign parity_check_matrix[0] = 11'b11111111111;
    assign parity_check_matrix[1] = 11'b00000000111;
    assign parity_check_matrix[2] = 11'b11111111001;
    assign parity_check_matrix[3] = 11'b00000001110;
    assign parity_check_matrix[4] = 11'b11111110000;
    assign parity_check_matrix[5] = 11'b00000001011;
    assign parity_check_matrix[6] = 11'b11111110101;
    assign parity_check_matrix[7] = 11'b00000010110;
    assign parity_check_matrix[8] = 11'b11111101000;
    assign parity_check_matrix[9] = 11'b00000010011;
    assign parity_check_matrix[10] = 11'b11111101101;
    assign parity_check_matrix[11] = 11'b00000100110;
    assign parity_check_matrix[12] = 11'b11111011000;
    assign parity_check_matrix[13] = 11'b00000100011;
    assign parity_check_matrix[14] = 11'b11111011101;
    assign parity_check_matrix[15] = 11'b00001000110;
    assign parity_check_matrix[16] = 11'b11110111000;
    assign parity_check_matrix[17] = 11'b00001000011;
    assign parity_check_matrix[18] = 11'b11110111101;
    assign parity_check_matrix[19] = 11'b00010000110;
    assign parity_check_matrix[20] = 11'b11101111000;
    assign parity_check_matrix[21] = 11'b00010000011;
    assign parity_check_matrix[22] = 11'b11101111101;
    assign parity_check_matrix[23] = 11'b00100000110;
    assign parity_check_matrix[24] = 11'b11011111000;
    assign parity_check_matrix[25] = 11'b00100000011;
    assign parity_check_matrix[26] = 11'b11011111101;
    assign parity_check_matrix[27] = 11'b01000000110;
    assign parity_check_matrix[28] = 11'b10111111000;
    assign parity_check_matrix[29] = 11'b01000000011;
    assign parity_check_matrix[30] = 11'b10111111101;
    assign parity_check_matrix[31] = 11'b10000000110;
    assign parity_check_matrix[32] = 11'b01111111000;
    assign parity_check_matrix[33] = 11'b10000000011;
    assign parity_check_matrix[34] = 11'b01111111101;
    assign parity_check_matrix[35] = 11'b00000011010;
    assign parity_check_matrix[36] = 11'b11111100100;
    assign parity_check_matrix[37] = 11'b00000001101;
    assign parity_check_matrix[38] = 11'b11111110011;
    assign parity_check_matrix[39] = 11'b00000101010;
    assign parity_check_matrix[40] = 11'b11111010100;
    assign parity_check_matrix[41] = 11'b00000010101;
    assign parity_check_matrix[42] = 11'b11111101011;
    assign parity_check_matrix[43] = 11'b00001001010;
    assign parity_check_matrix[44] = 11'b11110110100;
    assign parity_check_matrix[45] = 11'b00000100101;
    assign parity_check_matrix[46] = 11'b11111011011;
    assign parity_check_matrix[47] = 11'b00010001010;
    assign parity_check_matrix[48] = 11'b11101110100;
    assign parity_check_matrix[49] = 11'b00001000101;
    assign parity_check_matrix[50] = 11'b11110111011;
    assign parity_check_matrix[51] = 11'b00100001010;
    assign parity_check_matrix[52] = 11'b11011110100;
    assign parity_check_matrix[53] = 11'b00010000101;
    assign parity_check_matrix[54] = 11'b11101111011;
    assign parity_check_matrix[55] = 11'b01000001010;
    assign parity_check_matrix[56] = 11'b10111110100;
    assign parity_check_matrix[57] = 11'b00100000101;
    assign parity_check_matrix[58] = 11'b11011111011;
    assign parity_check_matrix[59] = 11'b10000001010;
    assign parity_check_matrix[60] = 11'b01111110100;
    assign parity_check_matrix[61] = 11'b01000000101;
    assign parity_check_matrix[62] = 11'b10111111011;
    assign parity_check_matrix[63] = 11'b00000110010;
    assign parity_check_matrix[64] = 11'b11111001100;
    assign parity_check_matrix[65] = 11'b10000000101;
    assign parity_check_matrix[66] = 11'b01111111011;
    assign parity_check_matrix[67] = 11'b00001010010;
    assign parity_check_matrix[68] = 11'b11110101100;
    assign parity_check_matrix[69] = 11'b00000011001;
    assign parity_check_matrix[70] = 11'b11111100111;
    assign parity_check_matrix[71] = 11'b00010010010;
    assign parity_check_matrix[72] = 11'b11101101100;
    assign parity_check_matrix[73] = 11'b00000101001;
    assign parity_check_matrix[74] = 11'b11111010111;
    assign parity_check_matrix[75] = 11'b00100010010;
    assign parity_check_matrix[76] = 11'b11011101100;
    assign parity_check_matrix[77] = 11'b00001001001;
    assign parity_check_matrix[78] = 11'b11110110111;
    assign parity_check_matrix[79] = 11'b01000010010;
    assign parity_check_matrix[80] = 11'b10111101100;
    assign parity_check_matrix[81] = 11'b00010001001;
    assign parity_check_matrix[82] = 11'b11101110111;
    assign parity_check_matrix[83] = 11'b10000010010;
    assign parity_check_matrix[84] = 11'b01111101100;
    assign parity_check_matrix[85] = 11'b00100001001;
    assign parity_check_matrix[86] = 11'b11011110111;
    assign parity_check_matrix[87] = 11'b00001100010;
    assign parity_check_matrix[88] = 11'b11110011100;
    assign parity_check_matrix[89] = 11'b01000001001;
    assign parity_check_matrix[90] = 11'b10111110111;
    assign parity_check_matrix[91] = 11'b00010100010;
    assign parity_check_matrix[92] = 11'b11101011100;
    assign parity_check_matrix[93] = 11'b10000001001;
    assign parity_check_matrix[94] = 11'b01111110111;
    assign parity_check_matrix[95] = 11'b00100100010;
    assign parity_check_matrix[96] = 11'b11011011100;
    assign parity_check_matrix[97] = 11'b00000110001;
    assign parity_check_matrix[98] = 11'b11111001111;
    assign parity_check_matrix[99] = 11'b01000100010;
    assign parity_check_matrix[100] = 11'b10111011100;
    assign parity_check_matrix[101] = 11'b00001010001;
    assign parity_check_matrix[102] = 11'b11110101111;
    assign parity_check_matrix[103] = 11'b10000100010;
    assign parity_check_matrix[104] = 11'b01111011100;
    assign parity_check_matrix[105] = 11'b00010010001;
    assign parity_check_matrix[106] = 11'b11101101111;
    assign parity_check_matrix[107] = 11'b00011000010;
    assign parity_check_matrix[108] = 11'b11100111100;
    assign parity_check_matrix[109] = 11'b00100010001;
    assign parity_check_matrix[110] = 11'b11011101111;
    assign parity_check_matrix[111] = 11'b00101000010;
    assign parity_check_matrix[112] = 11'b11010111100;
    assign parity_check_matrix[113] = 11'b01000010001;
    assign parity_check_matrix[114] = 11'b10111101111;
    assign parity_check_matrix[115] = 11'b01001000010;
    assign parity_check_matrix[116] = 11'b10110111100;
    assign parity_check_matrix[117] = 11'b10000010001;
    assign parity_check_matrix[118] = 11'b01111101111;
    assign parity_check_matrix[119] = 11'b10001000010;
    assign parity_check_matrix[120] = 11'b01110111100;
    assign parity_check_matrix[121] = 11'b00001100001;
    assign parity_check_matrix[122] = 11'b11110011111;
    assign parity_check_matrix[123] = 11'b00110000010;
    assign parity_check_matrix[124] = 11'b11001111100;
    assign parity_check_matrix[125] = 11'b00010100001;
    assign parity_check_matrix[126] = 11'b11101011111;
    assign parity_check_matrix[127] = 11'b01010000010;
    assign parity_check_matrix[128] = 11'b10101111100;
    assign parity_check_matrix[129] = 11'b00100100001;
    assign parity_check_matrix[130] = 11'b11011011111;
    assign parity_check_matrix[131] = 11'b10010000010;
    assign parity_check_matrix[132] = 11'b01101111100;
    assign parity_check_matrix[133] = 11'b01000100001;
    assign parity_check_matrix[134] = 11'b10111011111;
    assign parity_check_matrix[135] = 11'b01100000010;
    assign parity_check_matrix[136] = 11'b10011111100;
    assign parity_check_matrix[137] = 11'b10000100001;
    assign parity_check_matrix[138] = 11'b01111011111;
    assign parity_check_matrix[139] = 11'b10100000010;
    assign parity_check_matrix[140] = 11'b01011111100;
    assign parity_check_matrix[141] = 11'b00011000001;
    assign parity_check_matrix[142] = 11'b11100111111;
    assign parity_check_matrix[143] = 11'b11000000010;
    assign parity_check_matrix[144] = 11'b00111111100;
    assign parity_check_matrix[145] = 11'b00101000001;
    assign parity_check_matrix[146] = 11'b11010111111;
    assign parity_check_matrix[147] = 11'b00000011100;
    assign parity_check_matrix[148] = 11'b11111100010;
    assign parity_check_matrix[149] = 11'b01001000001;
    assign parity_check_matrix[150] = 11'b10110111111;
    assign parity_check_matrix[151] = 11'b00000101100;
    assign parity_check_matrix[152] = 11'b11111010010;
    assign parity_check_matrix[153] = 11'b10001000001;
    assign parity_check_matrix[154] = 11'b01110111111;
    assign parity_check_matrix[155] = 11'b00001001100;
    assign parity_check_matrix[156] = 11'b11110110010;
    assign parity_check_matrix[157] = 11'b00110000001;
    assign parity_check_matrix[158] = 11'b11001111111;
    assign parity_check_matrix[159] = 11'b00010001100;
    assign parity_check_matrix[160] = 11'b11101110010;
    assign parity_check_matrix[161] = 11'b01010000001;
    assign parity_check_matrix[162] = 11'b10101111111;
    assign parity_check_matrix[163] = 11'b00100001100;
    assign parity_check_matrix[164] = 11'b11011110010;
    assign parity_check_matrix[165] = 11'b10010000001;
    assign parity_check_matrix[166] = 11'b01101111111;
    assign parity_check_matrix[167] = 11'b01000001100;
    assign parity_check_matrix[168] = 11'b10111110010;
    assign parity_check_matrix[169] = 11'b01100000001;
    assign parity_check_matrix[170] = 11'b10011111111;
    assign parity_check_matrix[171] = 11'b10000001100;
    assign parity_check_matrix[172] = 11'b01111110010;
    assign parity_check_matrix[173] = 11'b10100000001;
    assign parity_check_matrix[174] = 11'b01011111111;
    assign parity_check_matrix[175] = 11'b00000110100;
    assign parity_check_matrix[176] = 11'b11111001010;
    assign parity_check_matrix[177] = 11'b11000000001;
    assign parity_check_matrix[178] = 11'b00111111111;
    assign parity_check_matrix[179] = 11'b00001010100;
    assign parity_check_matrix[180] = 11'b11110101010;
    assign parity_check_matrix[181] = 11'b00010010100;
    assign parity_check_matrix[182] = 11'b00001101000;
    assign parity_check_matrix[183] = 11'b11100000011;
    assign parity_check_matrix[184] = 11'b00100010100;
    assign parity_check_matrix[185] = 11'b00010101000;
    assign parity_check_matrix[186] = 11'b11001000011;
    assign parity_check_matrix[187] = 11'b01000010100;
    assign parity_check_matrix[188] = 11'b00100101000;
    assign parity_check_matrix[189] = 11'b10011000011;
    assign parity_check_matrix[190] = 11'b10000010100;
    assign parity_check_matrix[191] = 11'b01000101000;
    assign parity_check_matrix[192] = 11'b00111000011;
    assign parity_check_matrix[193] = 11'b00001100100;
    assign parity_check_matrix[194] = 11'b00010011000;
    assign parity_check_matrix[195] = 11'b11100001111;
    assign parity_check_matrix[196] = 11'b00001110000;
    assign parity_check_matrix[197] = 11'b11110000111;
    assign parity_check_matrix[198] = 11'b00000111000;
    assign parity_check_matrix[199] = 11'b11111000011;
    assign parity_check_matrix[200] = 11'b00010100100;
    assign parity_check_matrix[201] = 11'b00001011000;
    assign parity_check_matrix[202] = 11'b11100010111;
    assign parity_check_matrix[203] = 11'b10000101000;
    assign parity_check_matrix[204] = 11'b01111000111;
    assign parity_check_matrix[205] = 11'b00100011000;
    assign parity_check_matrix[206] = 11'b11011100011;
    assign parity_check_matrix[207] = 11'b00100100100;
    assign parity_check_matrix[208] = 11'b01000011000;
    assign parity_check_matrix[209] = 11'b10011001111;
    assign parity_check_matrix[210] = 11'b00010110000;
    assign parity_check_matrix[211] = 11'b11101000111;
    assign parity_check_matrix[212] = 11'b10000011000;
    assign parity_check_matrix[213] = 11'b01111100011;
    assign parity_check_matrix[214] = 11'b01000100100;
    assign parity_check_matrix[215] = 11'b00011001000;
    assign parity_check_matrix[216] = 11'b10100010011;
    assign parity_check_matrix[217] = 11'b10000100100;
    assign parity_check_matrix[218] = 11'b00101001000;
    assign parity_check_matrix[219] = 11'b01010010011;
    assign parity_check_matrix[220] = 11'b00011000100;
    assign parity_check_matrix[221] = 11'b01100001000;
    assign parity_check_matrix[222] = 11'b10000110011;
    assign parity_check_matrix[223] = 11'b00101000100;
    assign parity_check_matrix[224] = 11'b01010001000;
    assign parity_check_matrix[225] = 11'b10000111111;
    assign parity_check_matrix[226] = 11'b00100110000;
    assign parity_check_matrix[227] = 11'b11011000111;
    assign parity_check_matrix[228] = 11'b01001001000;
    assign parity_check_matrix[229] = 11'b10110110011;
    assign parity_check_matrix[230] = 11'b01001000100;
    assign parity_check_matrix[231] = 11'b00110001000;
    assign parity_check_matrix[232] = 11'b10001110111;
    assign parity_check_matrix[233] = 11'b10010001000;
    assign parity_check_matrix[234] = 11'b01100110111;
    assign parity_check_matrix[235] = 11'b10001001000;
    assign parity_check_matrix[236] = 11'b01110110011;
    assign parity_check_matrix[237] = 11'b10001000100;
    assign parity_check_matrix[238] = 11'b01000110000;
    assign parity_check_matrix[239] = 11'b00110001011;
    assign parity_check_matrix[240] = 11'b00110000100;
    assign parity_check_matrix[241] = 11'b11000001000;
    assign parity_check_matrix[242] = 11'b00001110011;
    assign parity_check_matrix[243] = 11'b01010000100;
    assign parity_check_matrix[244] = 11'b10100001000;
    assign parity_check_matrix[245] = 11'b00001111111;
    assign parity_check_matrix[246] = 11'b10000110000;
    assign parity_check_matrix[247] = 11'b01111001011;
    assign parity_check_matrix[248] = 11'b10010000100;
    assign parity_check_matrix[249] = 11'b01101110011;
    assign parity_check_matrix[250] = 11'b01100000100;
    assign parity_check_matrix[251] = 11'b00011010000;
    assign parity_check_matrix[252] = 11'b10000101011;
    assign parity_check_matrix[253] = 11'b10100000100;
    assign parity_check_matrix[254] = 11'b01001010000;
    assign parity_check_matrix[255] = 11'b00010101011;
    assign parity_check_matrix[256] = 11'b11000000100;
    assign parity_check_matrix[257] = 11'b00101010000;
    assign parity_check_matrix[258] = 11'b00010111111;
    assign parity_check_matrix[259] = 11'b00011100000;
    assign parity_check_matrix[260] = 11'b11100011011;
    assign parity_check_matrix[261] = 11'b00101100000;
    assign parity_check_matrix[262] = 11'b11010001111;
    assign parity_check_matrix[263] = 11'b10001010000;
    assign parity_check_matrix[264] = 11'b00110100000;
    assign parity_check_matrix[265] = 11'b01000001111;
    assign parity_check_matrix[266] = 11'b00110010000;
    assign parity_check_matrix[267] = 11'b01001100000;
    assign parity_check_matrix[268] = 11'b10000001111;
    assign parity_check_matrix[269] = 11'b01010010000;
    assign parity_check_matrix[270] = 11'b10001100000;
    assign parity_check_matrix[271] = 11'b00100001111;
    assign parity_check_matrix[272] = 11'b10010010000;
    assign parity_check_matrix[273] = 11'b01100100000;
    assign parity_check_matrix[274] = 11'b00001001111;
    assign parity_check_matrix[275] = 11'b01100010000;
    assign parity_check_matrix[276] = 11'b10010100000;
    assign parity_check_matrix[277] = 11'b00011011111;
    assign parity_check_matrix[278] = 11'b10100100000;
    assign parity_check_matrix[279] = 11'b01001011111;
    assign parity_check_matrix[280] = 11'b01010100000;
    assign parity_check_matrix[281] = 11'b10101001111;
    assign parity_check_matrix[282] = 11'b10100010000;
    assign parity_check_matrix[283] = 11'b01011000000;
    assign parity_check_matrix[284] = 11'b00000101111;
    assign parity_check_matrix[285] = 11'b11000010000;
    assign parity_check_matrix[286] = 11'b00111000000;
    assign parity_check_matrix[287] = 11'b00100111111;
    assign parity_check_matrix[288] = 11'b11000100000;
    assign parity_check_matrix[289] = 11'b00011101111;
    assign parity_check_matrix[290] = 11'b10011000000;
    assign parity_check_matrix[291] = 11'b01100011111;
    assign parity_check_matrix[292] = 11'b01101000000;
    assign parity_check_matrix[293] = 11'b00000011111;
    assign parity_check_matrix[294] = 11'b10010100011;
    assign parity_check_matrix[295] = 11'b11111111100;
    assign parity_check_matrix[296] = 11'b10101000000;
    assign parity_check_matrix[297] = 11'b00010001111;
    assign parity_check_matrix[298] = 11'b01000110011;
    assign parity_check_matrix[299] = 11'b11001000000;
    assign parity_check_matrix[300] = 11'b00110111101;
    assign parity_check_matrix[301] = 11'b01110000000;
    assign parity_check_matrix[302] = 11'b10001111110;
    assign parity_check_matrix[303] = 11'b10110000000;
    assign parity_check_matrix[304] = 11'b00000110111;
    assign parity_check_matrix[305] = 11'b01001001011;
    assign parity_check_matrix[306] = 11'b11010000000;
    assign parity_check_matrix[307] = 11'b00101111101;
    assign parity_check_matrix[308] = 11'b11100000000;
    assign parity_check_matrix[309] = 11'b00011111110;
    assign parity_check_matrix[310] = 11'b00001010111;
    assign parity_check_matrix[311] = 11'b11110101001;
    assign parity_check_matrix[312] = 11'b00000111110;
    assign parity_check_matrix[313] = 11'b11111000000;
    assign parity_check_matrix[314] = 11'b00010010111;
    assign parity_check_matrix[315] = 11'b11101101001;
    assign parity_check_matrix[316] = 11'b00001011110;
    assign parity_check_matrix[317] = 11'b11110100000;
    assign parity_check_matrix[318] = 11'b00100010111;
    assign parity_check_matrix[319] = 11'b11011101001;
    assign parity_check_matrix[320] = 11'b00010011110;
    assign parity_check_matrix[321] = 11'b11101100000;
    assign parity_check_matrix[322] = 11'b01000010111;
    assign parity_check_matrix[323] = 11'b10111101001;
    assign parity_check_matrix[324] = 11'b00100011110;
    assign parity_check_matrix[325] = 11'b11011100000;
    assign parity_check_matrix[326] = 11'b10000010111;
    assign parity_check_matrix[327] = 11'b01111101001;
    assign parity_check_matrix[328] = 11'b01000011110;
    assign parity_check_matrix[329] = 11'b10111100000;
    assign parity_check_matrix[330] = 11'b00001100111;
    assign parity_check_matrix[331] = 11'b11110011001;
    assign parity_check_matrix[332] = 11'b10000011110;
    assign parity_check_matrix[333] = 11'b01111100000;
    assign parity_check_matrix[334] = 11'b00010100111;
    assign parity_check_matrix[335] = 11'b11101011001;
    assign parity_check_matrix[336] = 11'b00001101110;
    assign parity_check_matrix[337] = 11'b11110010000;
    assign parity_check_matrix[338] = 11'b00100100111;
    assign parity_check_matrix[339] = 11'b11011011001;
    assign parity_check_matrix[340] = 11'b00010101110;
    assign parity_check_matrix[341] = 11'b11101010000;
    assign parity_check_matrix[342] = 11'b01000100111;
    assign parity_check_matrix[343] = 11'b10111011001;
    assign parity_check_matrix[344] = 11'b00100101110;
    assign parity_check_matrix[345] = 11'b11011010000;
    assign parity_check_matrix[346] = 11'b10000100111;
    assign parity_check_matrix[347] = 11'b01111011001;
    assign parity_check_matrix[348] = 11'b01000101110;
    assign parity_check_matrix[349] = 11'b10111010000;
    assign parity_check_matrix[350] = 11'b00011000111;
    assign parity_check_matrix[351] = 11'b11100111001;
    assign parity_check_matrix[352] = 11'b10000101110;
    assign parity_check_matrix[353] = 11'b01111010000;
    assign parity_check_matrix[354] = 11'b00101000111;
    assign parity_check_matrix[355] = 11'b11010111001;
    assign parity_check_matrix[356] = 11'b00011001110;
    assign parity_check_matrix[357] = 11'b11100110000;
    assign parity_check_matrix[358] = 11'b01001000111;
    assign parity_check_matrix[359] = 11'b10110111001;
    assign parity_check_matrix[360] = 11'b00101001110;
    assign parity_check_matrix[361] = 11'b11010110000;
    assign parity_check_matrix[362] = 11'b10001000111;
    assign parity_check_matrix[363] = 11'b01110111001;
    assign parity_check_matrix[364] = 11'b01001001110;
    assign parity_check_matrix[365] = 11'b10110110000;
    assign parity_check_matrix[366] = 11'b00110000111;
    assign parity_check_matrix[367] = 11'b11001111001;
    assign parity_check_matrix[368] = 11'b10001001110;
    assign parity_check_matrix[369] = 11'b01110110000;
    assign parity_check_matrix[370] = 11'b01010000111;
    assign parity_check_matrix[371] = 11'b10101111001;
    assign parity_check_matrix[372] = 11'b00110001110;
    assign parity_check_matrix[373] = 11'b11001110000;
    assign parity_check_matrix[374] = 11'b10010000111;
    assign parity_check_matrix[375] = 11'b01101111001;
    assign parity_check_matrix[376] = 11'b01010001110;
    assign parity_check_matrix[377] = 11'b10101110000;
    assign parity_check_matrix[378] = 11'b01100000111;
    assign parity_check_matrix[379] = 11'b10011111001;
    assign parity_check_matrix[380] = 11'b10010001110;
    assign parity_check_matrix[381] = 11'b01101110000;
    assign parity_check_matrix[382] = 11'b10100000111;
    assign parity_check_matrix[383] = 11'b01011111001;
    assign parity_check_matrix[384] = 11'b01100001110;
    assign parity_check_matrix[385] = 11'b10011110000;
    assign parity_check_matrix[386] = 11'b11000000111;
    assign parity_check_matrix[387] = 11'b00111111001;
    assign parity_check_matrix[388] = 11'b10100001110;
    assign parity_check_matrix[389] = 11'b01011110000;
    assign parity_check_matrix[390] = 11'b00000111011;
    assign parity_check_matrix[391] = 11'b11111000101;
    assign parity_check_matrix[392] = 11'b11000001110;
    assign parity_check_matrix[393] = 11'b00111110000;
    assign parity_check_matrix[394] = 11'b00001011011;
    assign parity_check_matrix[395] = 11'b11110100101;
    assign parity_check_matrix[396] = 11'b00001110110;
    assign parity_check_matrix[397] = 11'b11110001000;
    assign parity_check_matrix[398] = 11'b00010011011;
    assign parity_check_matrix[399] = 11'b11101100101;
    assign parity_check_matrix[400] = 11'b00010110110;
    assign parity_check_matrix[401] = 11'b11101001000;
    assign parity_check_matrix[402] = 11'b00100011011;
    assign parity_check_matrix[403] = 11'b11011100101;
    assign parity_check_matrix[404] = 11'b00100110110;
    assign parity_check_matrix[405] = 11'b11011001000;
    assign parity_check_matrix[406] = 11'b01000011011;
    assign parity_check_matrix[407] = 11'b10111100101;
    assign parity_check_matrix[408] = 11'b01000110110;
    assign parity_check_matrix[409] = 11'b10111001000;
    assign parity_check_matrix[410] = 11'b10000011011;
    assign parity_check_matrix[411] = 11'b01111100101;
    assign parity_check_matrix[412] = 11'b10000110110;
    assign parity_check_matrix[413] = 11'b01111001000;
    assign parity_check_matrix[414] = 11'b00001101011;
    assign parity_check_matrix[415] = 11'b11110010101;
    assign parity_check_matrix[416] = 11'b00011010110;
    assign parity_check_matrix[417] = 11'b11100101000;
    assign parity_check_matrix[418] = 11'b00100101011;
    assign parity_check_matrix[419] = 11'b11011010101;
    assign parity_check_matrix[420] = 11'b00101010110;
    assign parity_check_matrix[421] = 11'b11010101000;
    assign parity_check_matrix[422] = 11'b01000101011;
    assign parity_check_matrix[423] = 11'b10111010101;
    assign parity_check_matrix[424] = 11'b01001010110;
    assign parity_check_matrix[425] = 11'b10110101000;
    assign parity_check_matrix[426] = 11'b00011001011;
    assign parity_check_matrix[427] = 11'b11100110101;
    assign parity_check_matrix[428] = 11'b10001010110;
    assign parity_check_matrix[429] = 11'b01110101000;
    assign parity_check_matrix[430] = 11'b00101001011;
    assign parity_check_matrix[431] = 11'b11010110101;
    assign parity_check_matrix[432] = 11'b00110010110;
    assign parity_check_matrix[433] = 11'b11001101000;
    assign parity_check_matrix[434] = 11'b10001001011;
    assign parity_check_matrix[435] = 11'b01110110101;
    assign parity_check_matrix[436] = 11'b01010010110;
    assign parity_check_matrix[437] = 11'b10101101000;
    assign parity_check_matrix[438] = 11'b01010001011;
    assign parity_check_matrix[439] = 11'b10101110101;
    assign parity_check_matrix[440] = 11'b10010010110;
    assign parity_check_matrix[441] = 11'b01101101000;
    assign parity_check_matrix[442] = 11'b10010001011;
    assign parity_check_matrix[443] = 11'b01101110101;
    assign parity_check_matrix[444] = 11'b01100010110;
    assign parity_check_matrix[445] = 11'b10011101000;
    assign parity_check_matrix[446] = 11'b01100001011;
    assign parity_check_matrix[447] = 11'b10011110101;
    assign parity_check_matrix[448] = 11'b10100010110;
    assign parity_check_matrix[449] = 11'b01011101000;
    assign parity_check_matrix[450] = 11'b10100001011;
    assign parity_check_matrix[451] = 11'b01011110101;
    assign parity_check_matrix[452] = 11'b11000010110;
    assign parity_check_matrix[453] = 11'b00111101000;
    assign parity_check_matrix[454] = 11'b11000001011;
    assign parity_check_matrix[455] = 11'b00111110101;
    assign parity_check_matrix[456] = 11'b00011100110;
    assign parity_check_matrix[457] = 11'b11100011000;
    assign parity_check_matrix[458] = 11'b00010110011;
    assign parity_check_matrix[459] = 11'b11101001101;
    assign parity_check_matrix[460] = 11'b00101100110;
    assign parity_check_matrix[461] = 11'b11010011000;
    assign parity_check_matrix[462] = 11'b00100110011;
    assign parity_check_matrix[463] = 11'b11011001101;
    assign parity_check_matrix[464] = 11'b01001100110;
    assign parity_check_matrix[465] = 11'b10110011000;
    assign parity_check_matrix[466] = 11'b00011010011;
    assign parity_check_matrix[467] = 11'b11100101101;
    assign parity_check_matrix[468] = 11'b10001100110;
    assign parity_check_matrix[469] = 11'b01110011000;
    assign parity_check_matrix[470] = 11'b00101010011;
    assign parity_check_matrix[471] = 11'b11010101101;
    assign parity_check_matrix[472] = 11'b00110100110;
    assign parity_check_matrix[473] = 11'b11001011000;
    assign parity_check_matrix[474] = 11'b01001010011;
    assign parity_check_matrix[475] = 11'b10110101101;
    assign parity_check_matrix[476] = 11'b01010100110;
    assign parity_check_matrix[477] = 11'b10101011000;
    assign parity_check_matrix[478] = 11'b10001010011;
    assign parity_check_matrix[479] = 11'b01110101101;
    assign parity_check_matrix[480] = 11'b10010100110;
    assign parity_check_matrix[481] = 11'b01101011000;
    assign parity_check_matrix[482] = 11'b00110010011;
    assign parity_check_matrix[483] = 11'b11001101101;
    assign parity_check_matrix[484] = 11'b01100100110;
    assign parity_check_matrix[485] = 11'b10011011000;
    assign parity_check_matrix[486] = 11'b10010010011;
    assign parity_check_matrix[487] = 11'b01101101101;
    assign parity_check_matrix[488] = 11'b10100100110;
    assign parity_check_matrix[489] = 11'b01011011000;
    assign parity_check_matrix[490] = 11'b01100010011;
    assign parity_check_matrix[491] = 11'b10011101101;
    assign parity_check_matrix[492] = 11'b11000100110;
    assign parity_check_matrix[493] = 11'b00111011000;
    assign parity_check_matrix[494] = 11'b11000010011;
    assign parity_check_matrix[495] = 11'b00111101101;
    assign parity_check_matrix[496] = 11'b00111000110;
    assign parity_check_matrix[497] = 11'b11000111000;
    assign parity_check_matrix[498] = 11'b00011100011;
    assign parity_check_matrix[499] = 11'b11100011101;
    assign parity_check_matrix[500] = 11'b01011000110;
    assign parity_check_matrix[501] = 11'b10100111000;
    assign parity_check_matrix[502] = 11'b00101100011;
    assign parity_check_matrix[503] = 11'b11010011101;
    assign parity_check_matrix[504] = 11'b10011000110;
    assign parity_check_matrix[505] = 11'b01100111000;
    assign parity_check_matrix[506] = 11'b01001100011;
    assign parity_check_matrix[507] = 11'b10110011101;
    assign parity_check_matrix[508] = 11'b01101000110;
    assign parity_check_matrix[509] = 11'b10010111000;
    assign parity_check_matrix[510] = 11'b10001100011;
    assign parity_check_matrix[511] = 11'b01110011101;
    assign parity_check_matrix[512] = 11'b10101000110;
    assign parity_check_matrix[513] = 11'b01010111000;
    assign parity_check_matrix[514] = 11'b00110100011;
    assign parity_check_matrix[515] = 11'b11001011101;
    assign parity_check_matrix[516] = 11'b11001000110;
    assign parity_check_matrix[517] = 11'b00110111000;
    assign parity_check_matrix[518] = 11'b01010100011;
    assign parity_check_matrix[519] = 11'b10101011101;
    assign parity_check_matrix[520] = 11'b01110000110;
    assign parity_check_matrix[521] = 11'b10001111000;
    assign parity_check_matrix[522] = 11'b01100100011;
    assign parity_check_matrix[523] = 11'b10011011101;
    assign parity_check_matrix[524] = 11'b10110000110;
    assign parity_check_matrix[525] = 11'b01001111000;
    assign parity_check_matrix[526] = 11'b10100100011;
    assign parity_check_matrix[527] = 11'b01011011101;
    assign parity_check_matrix[528] = 11'b11010000110;
    assign parity_check_matrix[529] = 11'b00101111000;
    assign parity_check_matrix[530] = 11'b11000100011;
    assign parity_check_matrix[531] = 11'b00111011101;
    assign parity_check_matrix[532] = 11'b11100000110;
    assign parity_check_matrix[533] = 11'b00011111000;
    assign parity_check_matrix[534] = 11'b01011000011;
    assign parity_check_matrix[535] = 11'b10100111101;
    assign parity_check_matrix[536] = 11'b00001111010;
    assign parity_check_matrix[537] = 11'b11110000100;
    assign parity_check_matrix[538] = 11'b01101000011;
    assign parity_check_matrix[539] = 11'b10010111101;
    assign parity_check_matrix[540] = 11'b00010111010;
    assign parity_check_matrix[541] = 11'b11101000100;
    assign parity_check_matrix[542] = 11'b10101000011;
    assign parity_check_matrix[543] = 11'b01010111101;
    assign parity_check_matrix[544] = 11'b00100111010;
    assign parity_check_matrix[545] = 11'b11011000100;
    assign parity_check_matrix[546] = 11'b01110000011;
    assign parity_check_matrix[547] = 11'b10001111101;
    assign parity_check_matrix[548] = 11'b01000111010;
    assign parity_check_matrix[549] = 11'b10111000100;
    assign parity_check_matrix[550] = 11'b10110000011;
    assign parity_check_matrix[551] = 11'b01001111101;
    assign parity_check_matrix[552] = 11'b10000111010;
    assign parity_check_matrix[553] = 11'b01111000100;
    assign parity_check_matrix[554] = 11'b11010000011;
    assign parity_check_matrix[555] = 11'b00101111110;
    assign parity_check_matrix[556] = 11'b00000111101;
    assign parity_check_matrix[557] = 11'b11111001001;
    assign parity_check_matrix[558] = 11'b11111110110;
    assign parity_check_matrix[559] = 11'b00001011101;
    assign parity_check_matrix[560] = 11'b11110100011;
    assign parity_check_matrix[561] = 11'b00011011010;
    assign parity_check_matrix[562] = 11'b11100100100;
    assign parity_check_matrix[563] = 11'b00010011101;
    assign parity_check_matrix[564] = 11'b11101100011;
    assign parity_check_matrix[565] = 11'b00101011010;
    assign parity_check_matrix[566] = 11'b11010100100;
    assign parity_check_matrix[567] = 11'b00100011101;
    assign parity_check_matrix[568] = 11'b11011100110;
    assign parity_check_matrix[569] = 11'b00001111001;
    assign parity_check_matrix[570] = 11'b11110000010;
    assign parity_check_matrix[571] = 11'b01000011101;
    assign parity_check_matrix[572] = 11'b10111100011;
    assign parity_check_matrix[573] = 11'b01001011010;
    assign parity_check_matrix[574] = 11'b10110100100;
    assign parity_check_matrix[575] = 11'b10000011101;
    assign parity_check_matrix[576] = 11'b01111100110;
    assign parity_check_matrix[577] = 11'b00010111001;
    assign parity_check_matrix[578] = 11'b11101000010;
    assign parity_check_matrix[579] = 11'b00001101101;
    assign parity_check_matrix[580] = 11'b11110010011;
    assign parity_check_matrix[581] = 11'b10001011010;
    assign parity_check_matrix[582] = 11'b01110100100;
    assign parity_check_matrix[583] = 11'b00010101101;
    assign parity_check_matrix[584] = 11'b11101010011;
    assign parity_check_matrix[585] = 11'b00110011010;
    assign parity_check_matrix[586] = 11'b11001100100;
    assign parity_check_matrix[587] = 11'b00100101101;
    assign parity_check_matrix[588] = 11'b11011010011;
    assign parity_check_matrix[589] = 11'b01010011010;
    assign parity_check_matrix[590] = 11'b10101100100;
    assign parity_check_matrix[591] = 11'b01000101101;
    assign parity_check_matrix[592] = 11'b10111010011;
    assign parity_check_matrix[593] = 11'b10010011010;
    assign parity_check_matrix[594] = 11'b01101100100;
    assign parity_check_matrix[595] = 11'b10000101101;
    assign parity_check_matrix[596] = 11'b01111010011;
    assign parity_check_matrix[597] = 11'b01100011010;
    assign parity_check_matrix[598] = 11'b10011100100;
    assign parity_check_matrix[599] = 11'b00011001101;
    assign parity_check_matrix[600] = 11'b11100110011;
    assign parity_check_matrix[601] = 11'b10100011010;
    assign parity_check_matrix[602] = 11'b01011100100;
    assign parity_check_matrix[603] = 11'b00101001101;
    assign parity_check_matrix[604] = 11'b11010110011;
    assign parity_check_matrix[605] = 11'b11000011010;
    assign parity_check_matrix[606] = 11'b00111100100;
    assign parity_check_matrix[607] = 11'b01001001101;
    assign parity_check_matrix[608] = 11'b10110110110;
    assign parity_check_matrix[609] = 11'b00100111001;
    assign parity_check_matrix[610] = 11'b11011000010;
    assign parity_check_matrix[611] = 11'b10001001101;
    assign parity_check_matrix[612] = 11'b01110110110;
    assign parity_check_matrix[613] = 11'b01000111001;
    assign parity_check_matrix[614] = 11'b10111000010;
    assign parity_check_matrix[615] = 11'b00110001101;
    assign parity_check_matrix[616] = 11'b11001110011;
    assign parity_check_matrix[617] = 11'b00011101010;
    assign parity_check_matrix[618] = 11'b11100010100;
    assign parity_check_matrix[619] = 11'b01010001101;
    assign parity_check_matrix[620] = 11'b10101110011;
    assign parity_check_matrix[621] = 11'b00101101010;
    assign parity_check_matrix[622] = 11'b11010010100;
    assign parity_check_matrix[623] = 11'b10010001101;
    assign parity_check_matrix[624] = 11'b01101110110;
    assign parity_check_matrix[625] = 11'b10000111001;
    assign parity_check_matrix[626] = 11'b01111000010;
    assign parity_check_matrix[627] = 11'b01100001101;
    assign parity_check_matrix[628] = 11'b10011110011;
    assign parity_check_matrix[629] = 11'b01001101010;
    assign parity_check_matrix[630] = 11'b10110010100;
    assign parity_check_matrix[631] = 11'b10100001101;
    assign parity_check_matrix[632] = 11'b01011110011;
    assign parity_check_matrix[633] = 11'b10001101010;
    assign parity_check_matrix[634] = 11'b01110010100;
    assign parity_check_matrix[635] = 11'b11000001101;
    assign parity_check_matrix[636] = 11'b00111110011;
    assign parity_check_matrix[637] = 11'b00110101010;
    assign parity_check_matrix[638] = 11'b11001010100;
    assign parity_check_matrix[639] = 11'b00001110101;
    assign parity_check_matrix[640] = 11'b11110001011;
    assign parity_check_matrix[641] = 11'b01010101010;
    assign parity_check_matrix[642] = 11'b10101010100;
    assign parity_check_matrix[643] = 11'b00010110101;
    assign parity_check_matrix[644] = 11'b11101001011;
    assign parity_check_matrix[645] = 11'b10010101010;
    assign parity_check_matrix[646] = 11'b01101010100;
    assign parity_check_matrix[647] = 11'b00100110101;
    assign parity_check_matrix[648] = 11'b11011001011;
    assign parity_check_matrix[649] = 11'b01100101010;
    assign parity_check_matrix[650] = 11'b10011010100;
    assign parity_check_matrix[651] = 11'b01000110101;
    assign parity_check_matrix[652] = 11'b10111001011;
    assign parity_check_matrix[653] = 11'b10100101010;
    assign parity_check_matrix[654] = 11'b01011010100;
    assign parity_check_matrix[655] = 11'b10000110101;
    assign parity_check_matrix[656] = 11'b01111001110;
    assign parity_check_matrix[657] = 11'b00011011001;
    assign parity_check_matrix[658] = 11'b11100100010;
    assign parity_check_matrix[659] = 11'b00011010101;
    assign parity_check_matrix[660] = 11'b11100101011;
    assign parity_check_matrix[661] = 11'b11000101010;
    assign parity_check_matrix[662] = 11'b00111010100;
    assign parity_check_matrix[663] = 11'b00101010101;
    assign parity_check_matrix[664] = 11'b11010101011;
    assign parity_check_matrix[665] = 11'b00111001010;
    assign parity_check_matrix[666] = 11'b11000110100;
    assign parity_check_matrix[667] = 11'b01001010101;
    assign parity_check_matrix[668] = 11'b10110101011;
    assign parity_check_matrix[669] = 11'b01011001010;
    assign parity_check_matrix[670] = 11'b10100110100;
    assign parity_check_matrix[671] = 11'b10001010101;
    assign parity_check_matrix[672] = 11'b01110101011;
    assign parity_check_matrix[673] = 11'b10011001010;
    assign parity_check_matrix[674] = 11'b01100110100;
    assign parity_check_matrix[675] = 11'b00110010101;
    assign parity_check_matrix[676] = 11'b11001101011;
    assign parity_check_matrix[677] = 11'b01101001010;
    assign parity_check_matrix[678] = 11'b10010110100;
    assign parity_check_matrix[679] = 11'b01010010101;
    assign parity_check_matrix[680] = 11'b10101101011;
    assign parity_check_matrix[681] = 11'b10101001010;
    assign parity_check_matrix[682] = 11'b01010110100;
    assign parity_check_matrix[683] = 11'b10010010101;
    assign parity_check_matrix[684] = 11'b01101101011;
    assign parity_check_matrix[685] = 11'b11001001010;
    assign parity_check_matrix[686] = 11'b00110110100;
    assign parity_check_matrix[687] = 11'b01100010101;
    assign parity_check_matrix[688] = 11'b10011101011;
    assign parity_check_matrix[689] = 11'b01110001010;
    assign parity_check_matrix[690] = 11'b10001110100;
    assign parity_check_matrix[691] = 11'b10100010101;
    assign parity_check_matrix[692] = 11'b01011101011;
    assign parity_check_matrix[693] = 11'b10110001010;
    assign parity_check_matrix[694] = 11'b01001110100;
    assign parity_check_matrix[695] = 11'b11000010101;
    assign parity_check_matrix[696] = 11'b00111101011;
    assign parity_check_matrix[697] = 11'b11010001010;
    assign parity_check_matrix[698] = 11'b00101110100;
    assign parity_check_matrix[699] = 11'b00011100101;
    assign parity_check_matrix[700] = 11'b11100011110;
    assign parity_check_matrix[701] = 11'b00101011001;
    assign parity_check_matrix[702] = 11'b11010100010;
    assign parity_check_matrix[703] = 11'b00101100101;
    assign parity_check_matrix[704] = 11'b11010011011;
    assign parity_check_matrix[705] = 11'b11100001010;
    assign parity_check_matrix[706] = 11'b00011110100;
    assign parity_check_matrix[707] = 11'b01001100101;
    assign parity_check_matrix[708] = 11'b10110011011;
    assign parity_check_matrix[709] = 11'b00011110010;
    assign parity_check_matrix[710] = 11'b11100001100;
    assign parity_check_matrix[711] = 11'b10001100101;
    assign parity_check_matrix[712] = 11'b01110011011;
    assign parity_check_matrix[713] = 11'b00101110010;
    assign parity_check_matrix[714] = 11'b11010001100;
    assign parity_check_matrix[715] = 11'b00110100101;
    assign parity_check_matrix[716] = 11'b11001011011;
    assign parity_check_matrix[717] = 11'b01001110010;
    assign parity_check_matrix[718] = 11'b10110001100;
    assign parity_check_matrix[719] = 11'b01010100101;
    assign parity_check_matrix[720] = 11'b10101011011;
    assign parity_check_matrix[721] = 11'b10001110010;
    assign parity_check_matrix[722] = 11'b01110001100;
    assign parity_check_matrix[723] = 11'b10010100101;
    assign parity_check_matrix[724] = 11'b01101011011;
    assign parity_check_matrix[725] = 11'b00110110010;
    assign parity_check_matrix[726] = 11'b11001001100;
    assign parity_check_matrix[727] = 11'b01100100101;
    assign parity_check_matrix[728] = 11'b10011011011;
    assign parity_check_matrix[729] = 11'b01010110010;
    assign parity_check_matrix[730] = 11'b10101001100;
    assign parity_check_matrix[731] = 11'b10100100101;
    assign parity_check_matrix[732] = 11'b01011011011;
    assign parity_check_matrix[733] = 11'b10010110010;
    assign parity_check_matrix[734] = 11'b01101001100;
    assign parity_check_matrix[735] = 11'b11000100101;
    assign parity_check_matrix[736] = 11'b00111011011;
    assign parity_check_matrix[737] = 11'b01100110010;
    assign parity_check_matrix[738] = 11'b10011001100;
    assign parity_check_matrix[739] = 11'b00111000101;
    assign parity_check_matrix[740] = 11'b11000111011;
    assign parity_check_matrix[741] = 11'b10100110010;
    assign parity_check_matrix[742] = 11'b01011001100;
    assign parity_check_matrix[743] = 11'b01011000101;
    assign parity_check_matrix[744] = 11'b10100111011;
    assign parity_check_matrix[745] = 11'b11000110010;
    assign parity_check_matrix[746] = 11'b00111001100;
    assign parity_check_matrix[747] = 11'b10011000101;
    assign parity_check_matrix[748] = 11'b01100111011;
    assign parity_check_matrix[749] = 11'b00111010010;
    assign parity_check_matrix[750] = 11'b11000101100;
    assign parity_check_matrix[751] = 11'b01101000101;
    assign parity_check_matrix[752] = 11'b10010111011;
    assign parity_check_matrix[753] = 11'b01011010010;
    assign parity_check_matrix[754] = 11'b10100101100;
    assign parity_check_matrix[755] = 11'b10101000101;
    assign parity_check_matrix[756] = 11'b01010111011;
    assign parity_check_matrix[757] = 11'b10011010010;
    assign parity_check_matrix[758] = 11'b01100101100;
    assign parity_check_matrix[759] = 11'b11001000101;
    assign parity_check_matrix[760] = 11'b00110111011;
    assign parity_check_matrix[761] = 11'b01101010010;
    assign parity_check_matrix[762] = 11'b10010101100;
    assign parity_check_matrix[763] = 11'b01110000101;
    assign parity_check_matrix[764] = 11'b10001111011;
    assign parity_check_matrix[765] = 11'b10101010010;
    assign parity_check_matrix[766] = 11'b01010101100;
    assign parity_check_matrix[767] = 11'b10110000101;
    assign parity_check_matrix[768] = 11'b01001111011;
    assign parity_check_matrix[769] = 11'b11001010010;
    assign parity_check_matrix[770] = 11'b00110101100;
    assign parity_check_matrix[771] = 11'b11010000101;
    assign parity_check_matrix[772] = 11'b00101111011;
    assign parity_check_matrix[773] = 11'b01110010010;
    assign parity_check_matrix[774] = 11'b10001101100;
    assign parity_check_matrix[775] = 11'b11100000101;
    assign parity_check_matrix[776] = 11'b00011111011;
    assign parity_check_matrix[777] = 11'b10110010010;
    assign parity_check_matrix[778] = 11'b01001101100;
    assign parity_check_matrix[779] = 11'b01001011001;
    assign parity_check_matrix[780] = 11'b10110100111;
    assign parity_check_matrix[781] = 11'b11010010010;
    assign parity_check_matrix[782] = 11'b00101101100;
    assign parity_check_matrix[783] = 11'b10001011001;
    assign parity_check_matrix[784] = 11'b01110100111;
    assign parity_check_matrix[785] = 11'b11100010010;
    assign parity_check_matrix[786] = 11'b00011101100;
    assign parity_check_matrix[787] = 11'b00110011001;
    assign parity_check_matrix[788] = 11'b11001100111;
    assign parity_check_matrix[789] = 11'b00111100010;
    assign parity_check_matrix[790] = 11'b11000011100;
    assign parity_check_matrix[791] = 11'b01010011001;
    assign parity_check_matrix[792] = 11'b10101100111;
    assign parity_check_matrix[793] = 11'b01011100010;
    assign parity_check_matrix[794] = 11'b10100011100;
    assign parity_check_matrix[795] = 11'b10010011001;
    assign parity_check_matrix[796] = 11'b01101100111;
    assign parity_check_matrix[797] = 11'b10011100010;
    assign parity_check_matrix[798] = 11'b01100011100;
    assign parity_check_matrix[799] = 11'b01100011001;
    assign parity_check_matrix[800] = 11'b10011100111;
    assign parity_check_matrix[801] = 11'b01101100010;
    assign parity_check_matrix[802] = 11'b10010011100;
    assign parity_check_matrix[803] = 11'b10100011001;
    assign parity_check_matrix[804] = 11'b01011100111;
    assign parity_check_matrix[805] = 11'b10101100010;
    assign parity_check_matrix[806] = 11'b01010011100;
    assign parity_check_matrix[807] = 11'b11000011001;
    assign parity_check_matrix[808] = 11'b00111100111;
    assign parity_check_matrix[809] = 11'b11001100010;
    assign parity_check_matrix[810] = 11'b00110011100;
    assign parity_check_matrix[811] = 11'b00011101001;
    assign parity_check_matrix[812] = 11'b11100110110;
    assign parity_check_matrix[813] = 11'b00111001001;
    assign parity_check_matrix[814] = 11'b11000011111;
    assign parity_check_matrix[815] = 11'b01110100010;
    assign parity_check_matrix[816] = 11'b10001011100;
    assign parity_check_matrix[817] = 11'b00011110001;
    assign parity_check_matrix[818] = 11'b11100100111;
    assign parity_check_matrix[819] = 11'b11111011110;
    assign parity_check_matrix[820] = 11'b00101101001;
    assign parity_check_matrix[821] = 11'b11010010111;
    assign parity_check_matrix[822] = 11'b10110100010;
    assign parity_check_matrix[823] = 11'b01001011100;
    assign parity_check_matrix[824] = 11'b01001101001;
    assign parity_check_matrix[825] = 11'b10110010111;
    assign parity_check_matrix[826] = 11'b00001111100;
    assign parity_check_matrix[827] = 11'b11110001110;
    assign parity_check_matrix[828] = 11'b00101110001;
    assign parity_check_matrix[829] = 11'b11010100111;
    assign parity_check_matrix[830] = 11'b11111111010;
    assign parity_check_matrix[831] = 11'b01011001001;
    assign parity_check_matrix[832] = 11'b10100011111;
    assign parity_check_matrix[833] = 11'b00111110110;
    assign parity_check_matrix[834] = 11'b11000101001;
    assign parity_check_matrix[835] = 11'b01111010110;
    assign parity_check_matrix[836] = 11'b10001101001;
    assign parity_check_matrix[837] = 11'b11110010110;
    assign parity_check_matrix[838] = 11'b00110101001;
    assign parity_check_matrix[839] = 11'b11001010111;
    assign parity_check_matrix[840] = 11'b00010111100;
    assign parity_check_matrix[841] = 11'b11101001110;
    assign parity_check_matrix[842] = 11'b01001110001;
    assign parity_check_matrix[843] = 11'b10110001111;
    assign parity_check_matrix[844] = 11'b01010101001;
    assign parity_check_matrix[845] = 11'b10101110110;
    assign parity_check_matrix[846] = 11'b10010101001;
    assign parity_check_matrix[847] = 11'b11101010110;
    assign parity_check_matrix[848] = 11'b01111011010;
    assign parity_check_matrix[849] = 11'b10001110001;
    assign parity_check_matrix[850] = 11'b01110001111;
    assign parity_check_matrix[851] = 11'b01011110110;
    assign parity_check_matrix[852] = 11'b10100101001;
    assign parity_check_matrix[853] = 11'b10111010110;
    assign parity_check_matrix[854] = 11'b01100101001;
    assign parity_check_matrix[855] = 11'b11011010110;
    assign parity_check_matrix[856] = 11'b10011001001;
    assign parity_check_matrix[857] = 11'b01100111110;
    assign parity_check_matrix[858] = 11'b00110110001;
    assign parity_check_matrix[859] = 11'b11001001111;
    assign parity_check_matrix[860] = 11'b10011110110;
    assign parity_check_matrix[861] = 11'b01101001001;
    assign parity_check_matrix[862] = 11'b11110111110;
    assign parity_check_matrix[863] = 11'b01010110001;
    assign parity_check_matrix[864] = 11'b10101010111;
    assign parity_check_matrix[865] = 11'b11111101110;
    assign parity_check_matrix[866] = 11'b10101001001;
    assign parity_check_matrix[867] = 11'b01010110111;
    assign parity_check_matrix[868] = 11'b00100111100;
    assign parity_check_matrix[869] = 11'b11011001110;
    assign parity_check_matrix[870] = 11'b10010110001;
    assign parity_check_matrix[871] = 11'b01101001111;
    assign parity_check_matrix[872] = 11'b11001001001;
    assign parity_check_matrix[873] = 11'b00110110111;
    assign parity_check_matrix[874] = 11'b01000111100;
    assign parity_check_matrix[875] = 11'b10111000111;
    assign parity_check_matrix[876] = 11'b00111111010;
    assign parity_check_matrix[877] = 11'b11010001001;
    assign parity_check_matrix[878] = 11'b11101111110;
    assign parity_check_matrix[879] = 11'b01100110001;
    assign parity_check_matrix[880] = 11'b10111100110;
    assign parity_check_matrix[881] = 11'b11011011010;
    assign parity_check_matrix[882] = 11'b10100110001;
    assign parity_check_matrix[883] = 11'b01011001111;
    assign parity_check_matrix[884] = 11'b11001110110;
    assign parity_check_matrix[885] = 11'b01110001001;
    assign parity_check_matrix[886] = 11'b10111111110;
    assign parity_check_matrix[887] = 11'b11000110001;
    assign parity_check_matrix[888] = 11'b00111001111;
    assign parity_check_matrix[889] = 11'b11010110110;
    assign parity_check_matrix[890] = 11'b00111010001;
    assign parity_check_matrix[891] = 11'b01101101110;
    assign parity_check_matrix[892] = 11'b10110001001;
    assign parity_check_matrix[893] = 11'b11011111110;
    assign parity_check_matrix[894] = 11'b01101010001;
    assign parity_check_matrix[895] = 11'b10001101111;
    assign parity_check_matrix[896] = 11'b11110100110;
    assign parity_check_matrix[897] = 11'b01011010001;
    assign parity_check_matrix[898] = 11'b10100111110;
    assign parity_check_matrix[899] = 11'b11100001001;
    assign parity_check_matrix[900] = 11'b00011110111;
    assign parity_check_matrix[901] = 11'b10000111100;
    assign parity_check_matrix[902] = 11'b11111000110;
    assign parity_check_matrix[903] = 11'b01110010001;
    assign parity_check_matrix[904] = 11'b00101101111;
    assign parity_check_matrix[905] = 11'b01011111010;
    assign parity_check_matrix[906] = 11'b10011010001;
    assign parity_check_matrix[907] = 11'b11100101110;
    assign parity_check_matrix[908] = 11'b10101010001;
    assign parity_check_matrix[909] = 11'b01010101111;
    assign parity_check_matrix[910] = 11'b00011011100;
    assign parity_check_matrix[911] = 11'b11101100110;
    assign parity_check_matrix[912] = 11'b10110010001;
    assign parity_check_matrix[913] = 11'b01000111111;
    assign parity_check_matrix[914] = 11'b01111101010;
    assign parity_check_matrix[915] = 11'b11001010001;
    assign parity_check_matrix[916] = 11'b10110101110;
    assign parity_check_matrix[917] = 11'b11010010001;
    assign parity_check_matrix[918] = 11'b00111101110;
    assign parity_check_matrix[919] = 11'b11100010001;
    assign parity_check_matrix[920] = 11'b01001101111;
    assign parity_check_matrix[921] = 11'b00101011100;
    assign parity_check_matrix[922] = 11'b10010101111;
    assign parity_check_matrix[923] = 11'b00111100001;
    assign parity_check_matrix[924] = 11'b11000111110;
    assign parity_check_matrix[925] = 11'b01011100001;
    assign parity_check_matrix[926] = 11'b10101011110;
    assign parity_check_matrix[927] = 11'b11110011010;
    assign parity_check_matrix[928] = 11'b10011100001;
    assign parity_check_matrix[929] = 11'b01101010111;
    assign parity_check_matrix[930] = 11'b00110111110;
    assign parity_check_matrix[931] = 11'b11001100001;
    assign parity_check_matrix[932] = 11'b01110011110;
    assign parity_check_matrix[933] = 11'b10101100001;
    assign parity_check_matrix[934] = 11'b11010011110;
    assign parity_check_matrix[935] = 11'b01101100001;
    assign parity_check_matrix[936] = 11'b10010011111;
    assign parity_check_matrix[937] = 11'b01001111110;
    assign parity_check_matrix[938] = 11'b10110100001;
    assign parity_check_matrix[939] = 11'b00111011110;
    assign parity_check_matrix[940] = 11'b11010100001;
    assign parity_check_matrix[941] = 11'b01101011110;
    assign parity_check_matrix[942] = 11'b11100100001;
    assign parity_check_matrix[943] = 11'b10011011110;
    assign parity_check_matrix[944] = 11'b01110100001;
    assign parity_check_matrix[945] = 11'b10001011111;
    assign parity_check_matrix[946] = 11'b01010111110;
    assign parity_check_matrix[947] = 11'b10111000001;
    assign parity_check_matrix[948] = 11'b11001011110;
    assign parity_check_matrix[949] = 11'b00110101111;
    assign parity_check_matrix[950] = 11'b11101110001;
    assign parity_check_matrix[951] = 11'b10010111110;
    assign parity_check_matrix[952] = 11'b01111000001;
    assign parity_check_matrix[953] = 11'b10101101110;
    assign parity_check_matrix[954] = 11'b01010011111;
    assign parity_check_matrix[955] = 11'b11011000001;
    assign parity_check_matrix[956] = 11'b01101111010;
    assign parity_check_matrix[957] = 11'b10100110111;
    assign parity_check_matrix[958] = 11'b11101000001;
    assign parity_check_matrix[959] = 11'b01111111110;
    assign parity_check_matrix[960] = 11'b11110000001;
    assign parity_check_matrix[961] = 11'b00011111101;
    assign parity_check_matrix[962] = 11'b01011011110;
    assign parity_check_matrix[963] = 11'b10100101111;
    assign parity_check_matrix[964] = 11'b10011111010;
    assign parity_check_matrix[965] = 11'b00101011111;
    assign parity_check_matrix[966] = 11'b11000101111;
    assign parity_check_matrix[967] = 11'b11110110001;
    assign parity_check_matrix[968] = 11'b10110011110;
    assign parity_check_matrix[969] = 11'b01001110111;
    assign parity_check_matrix[970] = 11'b11111100001;
    assign parity_check_matrix[971] = 11'b01011101110;
    assign parity_check_matrix[972] = 11'b10110110101;
    assign parity_check_matrix[973] = 11'b11101011010;
    assign parity_check_matrix[974] = 11'b00110011111;
    assign parity_check_matrix[975] = 11'b11001110101;
    assign parity_check_matrix[976] = 11'b10011101110;
    assign parity_check_matrix[977] = 11'b01100101111;
    assign parity_check_matrix[978] = 11'b11111010001;
    assign parity_check_matrix[979] = 11'b11001101110;
    assign parity_check_matrix[980] = 11'b00111010111;
    assign parity_check_matrix[981] = 11'b00101110111;
    assign parity_check_matrix[982] = 11'b11110001101;
    assign parity_check_matrix[983] = 11'b11010111010;
    assign parity_check_matrix[984] = 11'b10010110111;
    assign parity_check_matrix[985] = 11'b01101011101;
    assign parity_check_matrix[986] = 11'b10101111010;
    assign parity_check_matrix[987] = 11'b01011010111;
    assign parity_check_matrix[988] = 11'b11000110111;
    assign parity_check_matrix[989] = 11'b01111001101;
    assign parity_check_matrix[990] = 11'b10110111010;
    assign parity_check_matrix[991] = 11'b10011010111;
    assign parity_check_matrix[992] = 11'b01100111101;
    assign parity_check_matrix[993] = 11'b11001111010;
    assign parity_check_matrix[994] = 11'b01110010111;
    assign parity_check_matrix[995] = 11'b10111101010;
    assign parity_check_matrix[996] = 11'b11000111101;
    assign parity_check_matrix[997] = 11'b10111001101;
    assign parity_check_matrix[998] = 11'b01111110001;
    assign parity_check_matrix[999] = 11'b01110101110;
    assign parity_check_matrix[1000] = 11'b10111011010;
    assign parity_check_matrix[1001] = 11'b11011110001;
    assign parity_check_matrix[1002] = 11'b11101101010;
    assign parity_check_matrix[1003] = 11'b01011101101;
    assign parity_check_matrix[1004] = 11'b10111001110;
    assign parity_check_matrix[1005] = 11'b11100111010;
    assign parity_check_matrix[1006] = 11'b10101101101;
    assign parity_check_matrix[1007] = 11'b01111010101;
    assign parity_check_matrix[1008] = 11'b11011101010;
    assign parity_check_matrix[1009] = 11'b11101010101;
    assign parity_check_matrix[1010] = 11'b01110111010;
    assign parity_check_matrix[1011] = 11'b10111110001;
    assign parity_check_matrix[1012] = 11'b11010101110;
    assign parity_check_matrix[1013] = 11'b10000000000;
    assign parity_check_matrix[1014] = 11'b01000000000;
    assign parity_check_matrix[1015] = 11'b00100000000;
    assign parity_check_matrix[1016] = 11'b00010000000;
    assign parity_check_matrix[1017] = 11'b00001000000;
    assign parity_check_matrix[1018] = 11'b00000100000;
    assign parity_check_matrix[1019] = 11'b00000010000;
    assign parity_check_matrix[1020] = 11'b00000001000;
    assign parity_check_matrix[1021] = 11'b00000000100;
    assign parity_check_matrix[1022] = 11'b00000000010;
    assign parity_check_matrix[1023] = 11'b00000000001;
  end else if ((CodewordWidth == 2048) && (MessageWidth == 2036)) begin : gen_2048_2036
    `BR_ASSERT_STATIC(parity_width_matches_a, ParityWidth == 12)
    assign syndrome[11] = cw[1] ^ cw[3] ^ cw[5] ^ cw[7] ^ cw[9] ^ cw[11] ^ cw[13] ^ cw[15] ^ cw[17] ^ cw[18] ^ cw[21] ^ cw[23] ^ cw[25] ^ cw[27] ^ cw[29] ^ cw[31] ^ cw[33] ^ cw[35] ^ cw[36] ^ cw[39] ^ cw[41] ^ cw[43] ^ cw[45] ^ cw[47] ^ cw[49] ^ cw[51] ^ cw[52] ^ cw[55] ^ cw[57] ^ cw[59] ^ cw[61] ^ cw[63] ^ cw[65] ^ cw[66] ^ cw[69] ^ cw[71] ^ cw[73] ^ cw[75] ^ cw[77] ^ cw[78] ^ cw[81] ^ cw[83] ^ cw[85] ^ cw[87] ^ cw[88] ^ cw[91] ^ cw[93] ^ cw[95] ^ cw[96] ^ cw[99] ^ cw[101] ^ cw[102] ^ cw[105] ^ cw[106] ^ cw[108] ^ cw[111] ^ cw[113] ^ cw[115] ^ cw[117] ^ cw[119] ^ cw[121] ^ cw[123] ^ cw[125] ^ cw[126] ^ cw[129] ^ cw[131] ^ cw[133] ^ cw[135] ^ cw[137] ^ cw[139] ^ cw[141] ^ cw[142] ^ cw[145] ^ cw[147] ^ cw[149] ^ cw[151] ^ cw[153] ^ cw[155] ^ cw[156] ^ cw[159] ^ cw[161] ^ cw[163] ^ cw[165] ^ cw[167] ^ cw[168] ^ cw[171] ^ cw[173] ^ cw[175] ^ cw[177] ^ cw[178] ^ cw[181] ^ cw[183] ^ cw[185] ^ cw[186] ^ cw[189] ^ cw[191] ^ cw[192] ^ cw[195] ^ cw[196] ^ cw[198] ^ cw[201] ^ cw[203] ^ cw[205] ^ cw[207] ^ cw[209] ^ cw[211] ^ cw[213] ^ cw[214] ^ cw[217] ^ cw[219] ^ cw[221] ^ cw[223] ^ cw[225] ^ cw[227] ^ cw[228] ^ cw[231] ^ cw[233] ^ cw[235] ^ cw[237] ^ cw[239] ^ cw[240] ^ cw[243] ^ cw[245] ^ cw[247] ^ cw[249] ^ cw[250] ^ cw[253] ^ cw[255] ^ cw[257] ^ cw[258] ^ cw[261] ^ cw[263] ^ cw[264] ^ cw[267] ^ cw[268] ^ cw[270] ^ cw[273] ^ cw[275] ^ cw[277] ^ cw[279] ^ cw[281] ^ cw[283] ^ cw[284] ^ cw[287] ^ cw[289] ^ cw[291] ^ cw[293] ^ cw[295] ^ cw[296] ^ cw[299] ^ cw[301] ^ cw[303] ^ cw[305] ^ cw[306] ^ cw[309] ^ cw[311] ^ cw[313] ^ cw[314] ^ cw[317] ^ cw[319] ^ cw[320] ^ cw[323] ^ cw[324] ^ cw[326] ^ cw[329] ^ cw[331] ^ cw[333] ^ cw[335] ^ cw[337] ^ cw[338] ^ cw[341] ^ cw[343] ^ cw[345] ^ cw[347] ^ cw[348] ^ cw[351] ^ cw[353] ^ cw[355] ^ cw[356] ^ cw[359] ^ cw[361] ^ cw[362] ^ cw[365] ^ cw[366] ^ cw[368] ^ cw[371] ^ cw[373] ^ cw[375] ^ cw[377] ^ cw[378] ^ cw[381] ^ cw[383] ^ cw[385] ^ cw[386] ^ cw[389] ^ cw[391] ^ cw[392] ^ cw[395] ^ cw[396] ^ cw[398] ^ cw[401] ^ cw[403] ^ cw[405] ^ cw[406] ^ cw[409] ^ cw[411] ^ cw[412] ^ cw[415] ^ cw[416] ^ cw[418] ^ cw[421] ^ cw[423] ^ cw[424] ^ cw[427] ^ cw[428] ^ cw[430] ^ cw[433] ^ cw[434] ^ cw[436] ^ cw[438] ^ cw[441] ^ cw[443] ^ cw[445] ^ cw[447] ^ cw[449] ^ cw[451] ^ cw[453] ^ cw[454] ^ cw[457] ^ cw[459] ^ cw[461] ^ cw[463] ^ cw[465] ^ cw[467] ^ cw[468] ^ cw[471] ^ cw[473] ^ cw[475] ^ cw[477] ^ cw[479] ^ cw[480] ^ cw[483] ^ cw[485] ^ cw[487] ^ cw[489] ^ cw[490] ^ cw[493] ^ cw[495] ^ cw[497] ^ cw[498] ^ cw[501] ^ cw[503] ^ cw[504] ^ cw[507] ^ cw[508] ^ cw[510] ^ cw[513] ^ cw[515] ^ cw[517] ^ cw[519] ^ cw[521] ^ cw[523] ^ cw[524] ^ cw[527] ^ cw[529] ^ cw[531] ^ cw[533] ^ cw[535] ^ cw[536] ^ cw[539] ^ cw[541] ^ cw[543] ^ cw[545] ^ cw[546] ^ cw[549] ^ cw[551] ^ cw[553] ^ cw[554] ^ cw[557] ^ cw[559] ^ cw[560] ^ cw[563] ^ cw[564] ^ cw[566] ^ cw[569] ^ cw[571] ^ cw[573] ^ cw[575] ^ cw[577] ^ cw[578] ^ cw[581] ^ cw[583] ^ cw[585] ^ cw[587] ^ cw[588] ^ cw[591] ^ cw[593] ^ cw[595] ^ cw[596] ^ cw[599] ^ cw[601] ^ cw[602] ^ cw[605] ^ cw[606] ^ cw[608] ^ cw[611] ^ cw[613] ^ cw[615] ^ cw[617] ^ cw[618] ^ cw[621] ^ cw[623] ^ cw[625] ^ cw[626] ^ cw[629] ^ cw[631] ^ cw[632] ^ cw[635] ^ cw[636] ^ cw[638] ^ cw[641] ^ cw[643] ^ cw[645] ^ cw[646] ^ cw[649] ^ cw[651] ^ cw[652] ^ cw[655] ^ cw[656] ^ cw[658] ^ cw[661] ^ cw[663] ^ cw[664] ^ cw[667] ^ cw[668] ^ cw[670] ^ cw[673] ^ cw[674] ^ cw[676] ^ cw[678] ^ cw[681] ^ cw[683] ^ cw[685] ^ cw[687] ^ cw[689] ^ cw[691] ^ cw[692] ^ cw[695] ^ cw[697] ^ cw[699] ^ cw[701] ^ cw[703] ^ cw[704] ^ cw[707] ^ cw[709] ^ cw[711] ^ cw[713] ^ cw[714] ^ cw[717] ^ cw[719] ^ cw[721] ^ cw[722] ^ cw[725] ^ cw[727] ^ cw[728] ^ cw[731] ^ cw[732] ^ cw[734] ^ cw[737] ^ cw[739] ^ cw[741] ^ cw[743] ^ cw[745] ^ cw[746] ^ cw[749] ^ cw[751] ^ cw[753] ^ cw[755] ^ cw[756] ^ cw[759] ^ cw[761] ^ cw[763] ^ cw[764] ^ cw[767] ^ cw[769] ^ cw[770] ^ cw[773] ^ cw[774] ^ cw[776] ^ cw[779] ^ cw[781] ^ cw[783] ^ cw[785] ^ cw[786] ^ cw[789] ^ cw[791] ^ cw[793] ^ cw[794] ^ cw[797] ^ cw[799] ^ cw[800] ^ cw[803] ^ cw[804] ^ cw[806] ^ cw[809] ^ cw[811] ^ cw[813] ^ cw[814] ^ cw[817] ^ cw[819] ^ cw[820] ^ cw[823] ^ cw[824] ^ cw[826] ^ cw[829] ^ cw[831] ^ cw[832] ^ cw[835] ^ cw[836] ^ cw[838] ^ cw[841] ^ cw[842] ^ cw[844] ^ cw[846] ^ cw[849] ^ cw[851] ^ cw[853] ^ cw[855] ^ cw[857] ^ cw[858] ^ cw[861] ^ cw[863] ^ cw[865] ^ cw[867] ^ cw[868] ^ cw[871] ^ cw[873] ^ cw[875] ^ cw[876] ^ cw[879] ^ cw[881] ^ cw[882] ^ cw[885] ^ cw[886] ^ cw[888] ^ cw[891] ^ cw[893] ^ cw[895] ^ cw[897] ^ cw[898] ^ cw[901] ^ cw[903] ^ cw[905] ^ cw[906] ^ cw[909] ^ cw[911] ^ cw[912] ^ cw[915] ^ cw[916] ^ cw[918] ^ cw[921] ^ cw[923] ^ cw[925] ^ cw[926] ^ cw[929] ^ cw[931] ^ cw[932] ^ cw[935] ^ cw[936] ^ cw[938] ^ cw[941] ^ cw[943] ^ cw[944] ^ cw[947] ^ cw[948] ^ cw[950] ^ cw[953] ^ cw[954] ^ cw[956] ^ cw[958] ^ cw[961] ^ cw[963] ^ cw[965] ^ cw[967] ^ cw[968] ^ cw[971] ^ cw[973] ^ cw[975] ^ cw[976] ^ cw[979] ^ cw[981] ^ cw[982] ^ cw[985] ^ cw[986] ^ cw[988] ^ cw[991] ^ cw[993] ^ cw[995] ^ cw[996] ^ cw[999] ^ cw[1001] ^ cw[1002] ^ cw[1005] ^ cw[1006] ^ cw[1008] ^ cw[1011] ^ cw[1013] ^ cw[1014] ^ cw[1017] ^ cw[1018] ^ cw[1020] ^ cw[1023] ^ cw[1024] ^ cw[1026] ^ cw[1028] ^ cw[1031] ^ cw[1033] ^ cw[1035] ^ cw[1036] ^ cw[1039] ^ cw[1041] ^ cw[1042] ^ cw[1045] ^ cw[1046] ^ cw[1048] ^ cw[1051] ^ cw[1053] ^ cw[1054] ^ cw[1057] ^ cw[1058] ^ cw[1060] ^ cw[1063] ^ cw[1064] ^ cw[1066] ^ cw[1068] ^ cw[1071] ^ cw[1073] ^ cw[1074] ^ cw[1077] ^ cw[1078] ^ cw[1080] ^ cw[1083] ^ cw[1084] ^ cw[1086] ^ cw[1088] ^ cw[1091] ^ cw[1092] ^ cw[1094] ^ cw[1096] ^ cw[1098] ^ cw[1101] ^ cw[1103] ^ cw[1105] ^ cw[1107] ^ cw[1109] ^ cw[1111] ^ cw[1112] ^ cw[1115] ^ cw[1117] ^ cw[1119] ^ cw[1121] ^ cw[1123] ^ cw[1124] ^ cw[1127] ^ cw[1129] ^ cw[1131] ^ cw[1133] ^ cw[1134] ^ cw[1137] ^ cw[1139] ^ cw[1141] ^ cw[1142] ^ cw[1145] ^ cw[1147] ^ cw[1148] ^ cw[1151] ^ cw[1152] ^ cw[1154] ^ cw[1157] ^ cw[1159] ^ cw[1161] ^ cw[1163] ^ cw[1165] ^ cw[1166] ^ cw[1169] ^ cw[1171] ^ cw[1173] ^ cw[1175] ^ cw[1176] ^ cw[1179] ^ cw[1181] ^ cw[1183] ^ cw[1184] ^ cw[1187] ^ cw[1189] ^ cw[1190] ^ cw[1193] ^ cw[1194] ^ cw[1196] ^ cw[1199] ^ cw[1201] ^ cw[1203] ^ cw[1205] ^ cw[1206] ^ cw[1209] ^ cw[1211] ^ cw[1213] ^ cw[1214] ^ cw[1217] ^ cw[1219] ^ cw[1220] ^ cw[1223] ^ cw[1224] ^ cw[1226] ^ cw[1229] ^ cw[1231] ^ cw[1233] ^ cw[1234] ^ cw[1237] ^ cw[1239] ^ cw[1240] ^ cw[1243] ^ cw[1244] ^ cw[1246] ^ cw[1249] ^ cw[1251] ^ cw[1252] ^ cw[1255] ^ cw[1256] ^ cw[1258] ^ cw[1261] ^ cw[1262] ^ cw[1264] ^ cw[1266] ^ cw[1269] ^ cw[1271] ^ cw[1273] ^ cw[1275] ^ cw[1277] ^ cw[1278] ^ cw[1281] ^ cw[1283] ^ cw[1285] ^ cw[1287] ^ cw[1288] ^ cw[1291] ^ cw[1293] ^ cw[1295] ^ cw[1296] ^ cw[1299] ^ cw[1301] ^ cw[1302] ^ cw[1305] ^ cw[1306] ^ cw[1308] ^ cw[1311] ^ cw[1313] ^ cw[1315] ^ cw[1317] ^ cw[1318] ^ cw[1321] ^ cw[1323] ^ cw[1325] ^ cw[1326] ^ cw[1329] ^ cw[1331] ^ cw[1332] ^ cw[1335] ^ cw[1336] ^ cw[1338] ^ cw[1341] ^ cw[1343] ^ cw[1345] ^ cw[1346] ^ cw[1349] ^ cw[1351] ^ cw[1352] ^ cw[1355] ^ cw[1356] ^ cw[1358] ^ cw[1361] ^ cw[1363] ^ cw[1364] ^ cw[1367] ^ cw[1368] ^ cw[1370] ^ cw[1373] ^ cw[1374] ^ cw[1376] ^ cw[1378] ^ cw[1381] ^ cw[1383] ^ cw[1385] ^ cw[1387] ^ cw[1388] ^ cw[1391] ^ cw[1393] ^ cw[1395] ^ cw[1396] ^ cw[1399] ^ cw[1401] ^ cw[1402] ^ cw[1405] ^ cw[1406] ^ cw[1408] ^ cw[1411] ^ cw[1413] ^ cw[1415] ^ cw[1416] ^ cw[1419] ^ cw[1421] ^ cw[1422] ^ cw[1425] ^ cw[1426] ^ cw[1428] ^ cw[1431] ^ cw[1433] ^ cw[1434] ^ cw[1437] ^ cw[1438] ^ cw[1440] ^ cw[1443] ^ cw[1444] ^ cw[1446] ^ cw[1448] ^ cw[1451] ^ cw[1453] ^ cw[1455] ^ cw[1456] ^ cw[1459] ^ cw[1461] ^ cw[1462] ^ cw[1465] ^ cw[1466] ^ cw[1468] ^ cw[1471] ^ cw[1473] ^ cw[1474] ^ cw[1477] ^ cw[1478] ^ cw[1480] ^ cw[1483] ^ cw[1484] ^ cw[1486] ^ cw[1488] ^ cw[1491] ^ cw[1493] ^ cw[1494] ^ cw[1497] ^ cw[1498] ^ cw[1500] ^ cw[1503] ^ cw[1504] ^ cw[1506] ^ cw[1508] ^ cw[1511] ^ cw[1512] ^ cw[1514] ^ cw[1516] ^ cw[1518] ^ cw[1521] ^ cw[1523] ^ cw[1525] ^ cw[1527] ^ cw[1529] ^ cw[1530] ^ cw[1533] ^ cw[1535] ^ cw[1537] ^ cw[1539] ^ cw[1540] ^ cw[1543] ^ cw[1545] ^ cw[1547] ^ cw[1548] ^ cw[1551] ^ cw[1553] ^ cw[1554] ^ cw[1557] ^ cw[1558] ^ cw[1560] ^ cw[1563] ^ cw[1565] ^ cw[1567] ^ cw[1569] ^ cw[1570] ^ cw[1573] ^ cw[1575] ^ cw[1577] ^ cw[1578] ^ cw[1581] ^ cw[1583] ^ cw[1584] ^ cw[1587] ^ cw[1588] ^ cw[1590] ^ cw[1593] ^ cw[1595] ^ cw[1597] ^ cw[1598] ^ cw[1601] ^ cw[1603] ^ cw[1604] ^ cw[1607] ^ cw[1608] ^ cw[1610] ^ cw[1613] ^ cw[1615] ^ cw[1616] ^ cw[1619] ^ cw[1620] ^ cw[1622] ^ cw[1625] ^ cw[1626] ^ cw[1628] ^ cw[1630] ^ cw[1633] ^ cw[1635] ^ cw[1637] ^ cw[1639] ^ cw[1640] ^ cw[1643] ^ cw[1645] ^ cw[1647] ^ cw[1648] ^ cw[1651] ^ cw[1653] ^ cw[1654] ^ cw[1657] ^ cw[1658] ^ cw[1660] ^ cw[1663] ^ cw[1665] ^ cw[1667] ^ cw[1668] ^ cw[1671] ^ cw[1673] ^ cw[1674] ^ cw[1677] ^ cw[1678] ^ cw[1680] ^ cw[1683] ^ cw[1685] ^ cw[1686] ^ cw[1689] ^ cw[1690] ^ cw[1692] ^ cw[1695] ^ cw[1696] ^ cw[1698] ^ cw[1700] ^ cw[1703] ^ cw[1705] ^ cw[1707] ^ cw[1708] ^ cw[1711] ^ cw[1713] ^ cw[1714] ^ cw[1717] ^ cw[1718] ^ cw[1720] ^ cw[1723] ^ cw[1725] ^ cw[1726] ^ cw[1729] ^ cw[1730] ^ cw[1732] ^ cw[1735] ^ cw[1736] ^ cw[1738] ^ cw[1740] ^ cw[1743] ^ cw[1745] ^ cw[1746] ^ cw[1749] ^ cw[1750] ^ cw[1752] ^ cw[1755] ^ cw[1756] ^ cw[1758] ^ cw[1760] ^ cw[1763] ^ cw[1764] ^ cw[1766] ^ cw[1768] ^ cw[1770] ^ cw[1773] ^ cw[1775] ^ cw[1777] ^ cw[1779] ^ cw[1780] ^ cw[1783] ^ cw[1785] ^ cw[1787] ^ cw[1788] ^ cw[1791] ^ cw[1793] ^ cw[1794] ^ cw[1797] ^ cw[1798] ^ cw[1800] ^ cw[1803] ^ cw[1805] ^ cw[1807] ^ cw[1808] ^ cw[1811] ^ cw[1813] ^ cw[1814] ^ cw[1817] ^ cw[1818] ^ cw[1820] ^ cw[1823] ^ cw[1825] ^ cw[1826] ^ cw[1829] ^ cw[1830] ^ cw[1832] ^ cw[1835] ^ cw[1836] ^ cw[1838] ^ cw[1840] ^ cw[1843] ^ cw[1845] ^ cw[1847] ^ cw[1848] ^ cw[1851] ^ cw[1853] ^ cw[1854] ^ cw[1857] ^ cw[1858] ^ cw[1860] ^ cw[1863] ^ cw[1865] ^ cw[1866] ^ cw[1869] ^ cw[1870] ^ cw[1872] ^ cw[1875] ^ cw[1876] ^ cw[1878] ^ cw[1880] ^ cw[1883] ^ cw[1885] ^ cw[1886] ^ cw[1889] ^ cw[1890] ^ cw[1892] ^ cw[1895] ^ cw[1896] ^ cw[1898] ^ cw[1900] ^ cw[1903] ^ cw[1904] ^ cw[1906] ^ cw[1908] ^ cw[1910] ^ cw[1913] ^ cw[1915] ^ cw[1917] ^ cw[1918] ^ cw[1921] ^ cw[1923] ^ cw[1924] ^ cw[1927] ^ cw[1928] ^ cw[1930] ^ cw[1933] ^ cw[1935] ^ cw[1936] ^ cw[1939] ^ cw[1940] ^ cw[1942] ^ cw[1945] ^ cw[1946] ^ cw[1948] ^ cw[1950] ^ cw[1953] ^ cw[1955] ^ cw[1956] ^ cw[1959] ^ cw[1960] ^ cw[1962] ^ cw[1965] ^ cw[1966] ^ cw[1968] ^ cw[1970] ^ cw[1973] ^ cw[1974] ^ cw[1976] ^ cw[1978] ^ cw[1980] ^ cw[1983] ^ cw[1985] ^ cw[1986] ^ cw[1989] ^ cw[1990] ^ cw[1992] ^ cw[1995] ^ cw[1996] ^ cw[1998] ^ cw[2000] ^ cw[2003] ^ cw[2004] ^ cw[2006] ^ cw[2008] ^ cw[2010] ^ cw[2013] ^ cw[2014] ^ cw[2016] ^ cw[2018] ^ cw[2020] ^ cw[2022] ^ cw[2025] ^ cw[2026] ^ cw[2027] ^ cw[2028] ^ cw[2029] ^ cw[2030] ^ cw[2031] ^ cw[2032] ^ cw[2033] ^ cw[2034] ^ cw[2035] ^ cw[2036];
    assign syndrome[10] = cw[1] ^ cw[3] ^ cw[5] ^ cw[7] ^ cw[9] ^ cw[11] ^ cw[13] ^ cw[15] ^ cw[16] ^ cw[19] ^ cw[21] ^ cw[23] ^ cw[25] ^ cw[27] ^ cw[29] ^ cw[31] ^ cw[33] ^ cw[34] ^ cw[37] ^ cw[39] ^ cw[41] ^ cw[43] ^ cw[45] ^ cw[47] ^ cw[49] ^ cw[50] ^ cw[53] ^ cw[55] ^ cw[57] ^ cw[59] ^ cw[61] ^ cw[63] ^ cw[64] ^ cw[67] ^ cw[69] ^ cw[71] ^ cw[73] ^ cw[75] ^ cw[76] ^ cw[79] ^ cw[81] ^ cw[83] ^ cw[85] ^ cw[86] ^ cw[89] ^ cw[91] ^ cw[93] ^ cw[94] ^ cw[97] ^ cw[99] ^ cw[100] ^ cw[103] ^ cw[104] ^ cw[107] ^ cw[108] ^ cw[111] ^ cw[113] ^ cw[115] ^ cw[117] ^ cw[119] ^ cw[121] ^ cw[123] ^ cw[124] ^ cw[127] ^ cw[129] ^ cw[131] ^ cw[133] ^ cw[135] ^ cw[137] ^ cw[139] ^ cw[140] ^ cw[143] ^ cw[145] ^ cw[147] ^ cw[149] ^ cw[151] ^ cw[153] ^ cw[154] ^ cw[157] ^ cw[159] ^ cw[161] ^ cw[163] ^ cw[165] ^ cw[166] ^ cw[169] ^ cw[171] ^ cw[173] ^ cw[175] ^ cw[176] ^ cw[179] ^ cw[181] ^ cw[183] ^ cw[184] ^ cw[187] ^ cw[189] ^ cw[190] ^ cw[193] ^ cw[194] ^ cw[197] ^ cw[198] ^ cw[201] ^ cw[203] ^ cw[205] ^ cw[207] ^ cw[209] ^ cw[211] ^ cw[212] ^ cw[215] ^ cw[217] ^ cw[219] ^ cw[221] ^ cw[223] ^ cw[225] ^ cw[226] ^ cw[229] ^ cw[231] ^ cw[233] ^ cw[235] ^ cw[237] ^ cw[238] ^ cw[241] ^ cw[243] ^ cw[245] ^ cw[247] ^ cw[248] ^ cw[251] ^ cw[253] ^ cw[255] ^ cw[256] ^ cw[259] ^ cw[261] ^ cw[262] ^ cw[265] ^ cw[266] ^ cw[269] ^ cw[270] ^ cw[273] ^ cw[275] ^ cw[277] ^ cw[279] ^ cw[281] ^ cw[282] ^ cw[285] ^ cw[287] ^ cw[289] ^ cw[291] ^ cw[293] ^ cw[294] ^ cw[297] ^ cw[299] ^ cw[301] ^ cw[303] ^ cw[304] ^ cw[307] ^ cw[309] ^ cw[311] ^ cw[312] ^ cw[315] ^ cw[317] ^ cw[318] ^ cw[321] ^ cw[322] ^ cw[325] ^ cw[326] ^ cw[329] ^ cw[331] ^ cw[333] ^ cw[335] ^ cw[336] ^ cw[339] ^ cw[341] ^ cw[343] ^ cw[345] ^ cw[346] ^ cw[349] ^ cw[351] ^ cw[353] ^ cw[354] ^ cw[357] ^ cw[359] ^ cw[360] ^ cw[363] ^ cw[364] ^ cw[367] ^ cw[368] ^ cw[371] ^ cw[373] ^ cw[375] ^ cw[376] ^ cw[379] ^ cw[381] ^ cw[383] ^ cw[384] ^ cw[387] ^ cw[389] ^ cw[390] ^ cw[393] ^ cw[394] ^ cw[397] ^ cw[398] ^ cw[401] ^ cw[403] ^ cw[404] ^ cw[407] ^ cw[409] ^ cw[410] ^ cw[413] ^ cw[414] ^ cw[417] ^ cw[418] ^ cw[421] ^ cw[422] ^ cw[425] ^ cw[426] ^ cw[429] ^ cw[430] ^ cw[432] ^ cw[435] ^ cw[436] ^ cw[438] ^ cw[441] ^ cw[443] ^ cw[445] ^ cw[447] ^ cw[449] ^ cw[451] ^ cw[452] ^ cw[455] ^ cw[457] ^ cw[459] ^ cw[461] ^ cw[463] ^ cw[465] ^ cw[466] ^ cw[469] ^ cw[471] ^ cw[473] ^ cw[475] ^ cw[477] ^ cw[478] ^ cw[481] ^ cw[483] ^ cw[485] ^ cw[487] ^ cw[488] ^ cw[491] ^ cw[493] ^ cw[495] ^ cw[496] ^ cw[499] ^ cw[501] ^ cw[502] ^ cw[505] ^ cw[506] ^ cw[509] ^ cw[510] ^ cw[513] ^ cw[515] ^ cw[517] ^ cw[519] ^ cw[521] ^ cw[522] ^ cw[525] ^ cw[527] ^ cw[529] ^ cw[531] ^ cw[533] ^ cw[534] ^ cw[537] ^ cw[539] ^ cw[541] ^ cw[543] ^ cw[544] ^ cw[547] ^ cw[549] ^ cw[551] ^ cw[552] ^ cw[555] ^ cw[557] ^ cw[558] ^ cw[561] ^ cw[562] ^ cw[565] ^ cw[566] ^ cw[569] ^ cw[571] ^ cw[573] ^ cw[575] ^ cw[576] ^ cw[579] ^ cw[581] ^ cw[583] ^ cw[585] ^ cw[586] ^ cw[589] ^ cw[591] ^ cw[593] ^ cw[594] ^ cw[597] ^ cw[599] ^ cw[600] ^ cw[603] ^ cw[604] ^ cw[607] ^ cw[608] ^ cw[611] ^ cw[613] ^ cw[615] ^ cw[616] ^ cw[619] ^ cw[621] ^ cw[623] ^ cw[624] ^ cw[627] ^ cw[629] ^ cw[630] ^ cw[633] ^ cw[634] ^ cw[637] ^ cw[638] ^ cw[641] ^ cw[643] ^ cw[644] ^ cw[647] ^ cw[649] ^ cw[650] ^ cw[653] ^ cw[654] ^ cw[657] ^ cw[658] ^ cw[661] ^ cw[662] ^ cw[665] ^ cw[666] ^ cw[669] ^ cw[670] ^ cw[672] ^ cw[675] ^ cw[676] ^ cw[678] ^ cw[681] ^ cw[683] ^ cw[685] ^ cw[687] ^ cw[689] ^ cw[690] ^ cw[693] ^ cw[695] ^ cw[697] ^ cw[699] ^ cw[701] ^ cw[702] ^ cw[705] ^ cw[707] ^ cw[709] ^ cw[711] ^ cw[712] ^ cw[715] ^ cw[717] ^ cw[719] ^ cw[720] ^ cw[723] ^ cw[725] ^ cw[726] ^ cw[729] ^ cw[730] ^ cw[733] ^ cw[734] ^ cw[737] ^ cw[739] ^ cw[741] ^ cw[743] ^ cw[744] ^ cw[747] ^ cw[749] ^ cw[751] ^ cw[753] ^ cw[754] ^ cw[757] ^ cw[759] ^ cw[761] ^ cw[762] ^ cw[765] ^ cw[767] ^ cw[768] ^ cw[771] ^ cw[772] ^ cw[775] ^ cw[776] ^ cw[779] ^ cw[781] ^ cw[783] ^ cw[784] ^ cw[787] ^ cw[789] ^ cw[791] ^ cw[792] ^ cw[795] ^ cw[797] ^ cw[798] ^ cw[801] ^ cw[802] ^ cw[805] ^ cw[806] ^ cw[809] ^ cw[811] ^ cw[812] ^ cw[815] ^ cw[817] ^ cw[818] ^ cw[821] ^ cw[822] ^ cw[825] ^ cw[826] ^ cw[829] ^ cw[830] ^ cw[833] ^ cw[834] ^ cw[837] ^ cw[838] ^ cw[840] ^ cw[843] ^ cw[844] ^ cw[846] ^ cw[849] ^ cw[851] ^ cw[853] ^ cw[855] ^ cw[856] ^ cw[859] ^ cw[861] ^ cw[863] ^ cw[865] ^ cw[866] ^ cw[869] ^ cw[871] ^ cw[873] ^ cw[874] ^ cw[877] ^ cw[879] ^ cw[880] ^ cw[883] ^ cw[884] ^ cw[887] ^ cw[888] ^ cw[891] ^ cw[893] ^ cw[895] ^ cw[896] ^ cw[899] ^ cw[901] ^ cw[903] ^ cw[904] ^ cw[907] ^ cw[909] ^ cw[910] ^ cw[913] ^ cw[914] ^ cw[917] ^ cw[918] ^ cw[921] ^ cw[923] ^ cw[924] ^ cw[927] ^ cw[929] ^ cw[930] ^ cw[933] ^ cw[934] ^ cw[937] ^ cw[938] ^ cw[941] ^ cw[942] ^ cw[945] ^ cw[946] ^ cw[949] ^ cw[950] ^ cw[952] ^ cw[955] ^ cw[956] ^ cw[958] ^ cw[961] ^ cw[963] ^ cw[965] ^ cw[966] ^ cw[969] ^ cw[971] ^ cw[973] ^ cw[974] ^ cw[977] ^ cw[979] ^ cw[980] ^ cw[983] ^ cw[984] ^ cw[987] ^ cw[988] ^ cw[991] ^ cw[993] ^ cw[994] ^ cw[997] ^ cw[999] ^ cw[1000] ^ cw[1003] ^ cw[1004] ^ cw[1007] ^ cw[1008] ^ cw[1011] ^ cw[1012] ^ cw[1015] ^ cw[1016] ^ cw[1019] ^ cw[1020] ^ cw[1022] ^ cw[1025] ^ cw[1026] ^ cw[1028] ^ cw[1031] ^ cw[1033] ^ cw[1034] ^ cw[1037] ^ cw[1039] ^ cw[1040] ^ cw[1043] ^ cw[1044] ^ cw[1047] ^ cw[1048] ^ cw[1051] ^ cw[1052] ^ cw[1055] ^ cw[1056] ^ cw[1059] ^ cw[1060] ^ cw[1062] ^ cw[1065] ^ cw[1066] ^ cw[1068] ^ cw[1071] ^ cw[1072] ^ cw[1075] ^ cw[1076] ^ cw[1079] ^ cw[1080] ^ cw[1082] ^ cw[1085] ^ cw[1086] ^ cw[1088] ^ cw[1090] ^ cw[1093] ^ cw[1094] ^ cw[1096] ^ cw[1098] ^ cw[1101] ^ cw[1103] ^ cw[1105] ^ cw[1107] ^ cw[1109] ^ cw[1110] ^ cw[1113] ^ cw[1115] ^ cw[1117] ^ cw[1119] ^ cw[1121] ^ cw[1122] ^ cw[1125] ^ cw[1127] ^ cw[1129] ^ cw[1131] ^ cw[1132] ^ cw[1135] ^ cw[1137] ^ cw[1139] ^ cw[1140] ^ cw[1143] ^ cw[1145] ^ cw[1146] ^ cw[1149] ^ cw[1150] ^ cw[1153] ^ cw[1154] ^ cw[1157] ^ cw[1159] ^ cw[1161] ^ cw[1163] ^ cw[1164] ^ cw[1167] ^ cw[1169] ^ cw[1171] ^ cw[1173] ^ cw[1174] ^ cw[1177] ^ cw[1179] ^ cw[1181] ^ cw[1182] ^ cw[1185] ^ cw[1187] ^ cw[1188] ^ cw[1191] ^ cw[1192] ^ cw[1195] ^ cw[1196] ^ cw[1199] ^ cw[1201] ^ cw[1203] ^ cw[1204] ^ cw[1207] ^ cw[1209] ^ cw[1211] ^ cw[1212] ^ cw[1215] ^ cw[1217] ^ cw[1218] ^ cw[1221] ^ cw[1222] ^ cw[1225] ^ cw[1226] ^ cw[1229] ^ cw[1231] ^ cw[1232] ^ cw[1235] ^ cw[1237] ^ cw[1238] ^ cw[1241] ^ cw[1242] ^ cw[1245] ^ cw[1246] ^ cw[1249] ^ cw[1250] ^ cw[1253] ^ cw[1254] ^ cw[1257] ^ cw[1258] ^ cw[1260] ^ cw[1263] ^ cw[1264] ^ cw[1266] ^ cw[1269] ^ cw[1271] ^ cw[1273] ^ cw[1275] ^ cw[1276] ^ cw[1279] ^ cw[1281] ^ cw[1283] ^ cw[1285] ^ cw[1286] ^ cw[1289] ^ cw[1291] ^ cw[1293] ^ cw[1294] ^ cw[1297] ^ cw[1299] ^ cw[1300] ^ cw[1303] ^ cw[1304] ^ cw[1307] ^ cw[1308] ^ cw[1311] ^ cw[1313] ^ cw[1315] ^ cw[1316] ^ cw[1319] ^ cw[1321] ^ cw[1323] ^ cw[1324] ^ cw[1327] ^ cw[1329] ^ cw[1330] ^ cw[1333] ^ cw[1334] ^ cw[1337] ^ cw[1338] ^ cw[1341] ^ cw[1343] ^ cw[1344] ^ cw[1347] ^ cw[1349] ^ cw[1350] ^ cw[1353] ^ cw[1354] ^ cw[1357] ^ cw[1358] ^ cw[1361] ^ cw[1362] ^ cw[1365] ^ cw[1366] ^ cw[1369] ^ cw[1370] ^ cw[1372] ^ cw[1375] ^ cw[1376] ^ cw[1378] ^ cw[1381] ^ cw[1383] ^ cw[1385] ^ cw[1386] ^ cw[1389] ^ cw[1391] ^ cw[1393] ^ cw[1394] ^ cw[1397] ^ cw[1399] ^ cw[1400] ^ cw[1403] ^ cw[1404] ^ cw[1407] ^ cw[1408] ^ cw[1411] ^ cw[1413] ^ cw[1414] ^ cw[1417] ^ cw[1419] ^ cw[1420] ^ cw[1423] ^ cw[1424] ^ cw[1427] ^ cw[1428] ^ cw[1431] ^ cw[1432] ^ cw[1435] ^ cw[1436] ^ cw[1439] ^ cw[1440] ^ cw[1442] ^ cw[1445] ^ cw[1446] ^ cw[1448] ^ cw[1451] ^ cw[1453] ^ cw[1454] ^ cw[1457] ^ cw[1459] ^ cw[1460] ^ cw[1463] ^ cw[1464] ^ cw[1467] ^ cw[1468] ^ cw[1471] ^ cw[1472] ^ cw[1475] ^ cw[1476] ^ cw[1479] ^ cw[1480] ^ cw[1482] ^ cw[1485] ^ cw[1486] ^ cw[1488] ^ cw[1491] ^ cw[1492] ^ cw[1495] ^ cw[1496] ^ cw[1499] ^ cw[1500] ^ cw[1502] ^ cw[1505] ^ cw[1506] ^ cw[1508] ^ cw[1510] ^ cw[1513] ^ cw[1514] ^ cw[1516] ^ cw[1518] ^ cw[1521] ^ cw[1523] ^ cw[1525] ^ cw[1527] ^ cw[1528] ^ cw[1531] ^ cw[1533] ^ cw[1535] ^ cw[1537] ^ cw[1538] ^ cw[1541] ^ cw[1543] ^ cw[1545] ^ cw[1546] ^ cw[1549] ^ cw[1551] ^ cw[1552] ^ cw[1555] ^ cw[1556] ^ cw[1559] ^ cw[1560] ^ cw[1563] ^ cw[1565] ^ cw[1567] ^ cw[1568] ^ cw[1571] ^ cw[1573] ^ cw[1575] ^ cw[1576] ^ cw[1579] ^ cw[1581] ^ cw[1582] ^ cw[1585] ^ cw[1586] ^ cw[1589] ^ cw[1590] ^ cw[1593] ^ cw[1595] ^ cw[1596] ^ cw[1599] ^ cw[1601] ^ cw[1602] ^ cw[1605] ^ cw[1606] ^ cw[1609] ^ cw[1610] ^ cw[1613] ^ cw[1614] ^ cw[1617] ^ cw[1618] ^ cw[1621] ^ cw[1622] ^ cw[1624] ^ cw[1627] ^ cw[1628] ^ cw[1630] ^ cw[1633] ^ cw[1635] ^ cw[1637] ^ cw[1638] ^ cw[1641] ^ cw[1643] ^ cw[1645] ^ cw[1646] ^ cw[1649] ^ cw[1651] ^ cw[1652] ^ cw[1655] ^ cw[1656] ^ cw[1659] ^ cw[1660] ^ cw[1663] ^ cw[1665] ^ cw[1666] ^ cw[1669] ^ cw[1671] ^ cw[1672] ^ cw[1675] ^ cw[1676] ^ cw[1679] ^ cw[1680] ^ cw[1683] ^ cw[1684] ^ cw[1687] ^ cw[1688] ^ cw[1691] ^ cw[1692] ^ cw[1694] ^ cw[1697] ^ cw[1698] ^ cw[1700] ^ cw[1703] ^ cw[1705] ^ cw[1706] ^ cw[1709] ^ cw[1711] ^ cw[1712] ^ cw[1715] ^ cw[1716] ^ cw[1719] ^ cw[1720] ^ cw[1723] ^ cw[1724] ^ cw[1727] ^ cw[1728] ^ cw[1731] ^ cw[1732] ^ cw[1734] ^ cw[1737] ^ cw[1738] ^ cw[1740] ^ cw[1743] ^ cw[1744] ^ cw[1747] ^ cw[1748] ^ cw[1751] ^ cw[1752] ^ cw[1754] ^ cw[1757] ^ cw[1758] ^ cw[1760] ^ cw[1762] ^ cw[1765] ^ cw[1766] ^ cw[1768] ^ cw[1770] ^ cw[1773] ^ cw[1775] ^ cw[1777] ^ cw[1778] ^ cw[1781] ^ cw[1783] ^ cw[1785] ^ cw[1786] ^ cw[1789] ^ cw[1791] ^ cw[1792] ^ cw[1795] ^ cw[1796] ^ cw[1799] ^ cw[1800] ^ cw[1803] ^ cw[1805] ^ cw[1806] ^ cw[1809] ^ cw[1811] ^ cw[1812] ^ cw[1815] ^ cw[1816] ^ cw[1819] ^ cw[1820] ^ cw[1823] ^ cw[1824] ^ cw[1827] ^ cw[1828] ^ cw[1831] ^ cw[1832] ^ cw[1834] ^ cw[1837] ^ cw[1838] ^ cw[1840] ^ cw[1843] ^ cw[1845] ^ cw[1846] ^ cw[1849] ^ cw[1851] ^ cw[1852] ^ cw[1855] ^ cw[1856] ^ cw[1859] ^ cw[1860] ^ cw[1863] ^ cw[1864] ^ cw[1867] ^ cw[1868] ^ cw[1871] ^ cw[1872] ^ cw[1874] ^ cw[1877] ^ cw[1878] ^ cw[1880] ^ cw[1883] ^ cw[1884] ^ cw[1887] ^ cw[1888] ^ cw[1891] ^ cw[1892] ^ cw[1894] ^ cw[1897] ^ cw[1898] ^ cw[1900] ^ cw[1902] ^ cw[1905] ^ cw[1906] ^ cw[1908] ^ cw[1910] ^ cw[1913] ^ cw[1915] ^ cw[1916] ^ cw[1919] ^ cw[1921] ^ cw[1922] ^ cw[1925] ^ cw[1926] ^ cw[1929] ^ cw[1930] ^ cw[1933] ^ cw[1934] ^ cw[1937] ^ cw[1938] ^ cw[1941] ^ cw[1942] ^ cw[1944] ^ cw[1947] ^ cw[1948] ^ cw[1950] ^ cw[1953] ^ cw[1954] ^ cw[1957] ^ cw[1958] ^ cw[1961] ^ cw[1962] ^ cw[1964] ^ cw[1967] ^ cw[1968] ^ cw[1970] ^ cw[1972] ^ cw[1975] ^ cw[1976] ^ cw[1978] ^ cw[1980] ^ cw[1983] ^ cw[1984] ^ cw[1987] ^ cw[1988] ^ cw[1991] ^ cw[1992] ^ cw[1994] ^ cw[1997] ^ cw[1998] ^ cw[2000] ^ cw[2002] ^ cw[2005] ^ cw[2006] ^ cw[2008] ^ cw[2010] ^ cw[2012] ^ cw[2015] ^ cw[2016] ^ cw[2018] ^ cw[2020] ^ cw[2022] ^ cw[2024] ^ cw[2026] ^ cw[2027] ^ cw[2028] ^ cw[2029] ^ cw[2030] ^ cw[2031] ^ cw[2032] ^ cw[2033] ^ cw[2034] ^ cw[2035] ^ cw[2037];
    assign syndrome[9] = cw[1] ^ cw[3] ^ cw[5] ^ cw[7] ^ cw[9] ^ cw[11] ^ cw[13] ^ cw[14] ^ cw[17] ^ cw[19] ^ cw[21] ^ cw[23] ^ cw[25] ^ cw[27] ^ cw[29] ^ cw[31] ^ cw[32] ^ cw[35] ^ cw[37] ^ cw[39] ^ cw[41] ^ cw[43] ^ cw[45] ^ cw[47] ^ cw[48] ^ cw[51] ^ cw[53] ^ cw[55] ^ cw[57] ^ cw[59] ^ cw[61] ^ cw[62] ^ cw[65] ^ cw[67] ^ cw[69] ^ cw[71] ^ cw[73] ^ cw[74] ^ cw[77] ^ cw[79] ^ cw[81] ^ cw[83] ^ cw[84] ^ cw[87] ^ cw[89] ^ cw[91] ^ cw[92] ^ cw[95] ^ cw[97] ^ cw[98] ^ cw[101] ^ cw[103] ^ cw[104] ^ cw[106] ^ cw[109] ^ cw[111] ^ cw[113] ^ cw[115] ^ cw[117] ^ cw[119] ^ cw[121] ^ cw[122] ^ cw[125] ^ cw[127] ^ cw[129] ^ cw[131] ^ cw[133] ^ cw[135] ^ cw[137] ^ cw[138] ^ cw[141] ^ cw[143] ^ cw[145] ^ cw[147] ^ cw[149] ^ cw[151] ^ cw[152] ^ cw[155] ^ cw[157] ^ cw[159] ^ cw[161] ^ cw[163] ^ cw[164] ^ cw[167] ^ cw[169] ^ cw[171] ^ cw[173] ^ cw[174] ^ cw[177] ^ cw[179] ^ cw[181] ^ cw[182] ^ cw[185] ^ cw[187] ^ cw[188] ^ cw[191] ^ cw[193] ^ cw[194] ^ cw[196] ^ cw[199] ^ cw[201] ^ cw[203] ^ cw[205] ^ cw[207] ^ cw[209] ^ cw[210] ^ cw[213] ^ cw[215] ^ cw[217] ^ cw[219] ^ cw[221] ^ cw[223] ^ cw[224] ^ cw[227] ^ cw[229] ^ cw[231] ^ cw[233] ^ cw[235] ^ cw[236] ^ cw[239] ^ cw[241] ^ cw[243] ^ cw[245] ^ cw[246] ^ cw[249] ^ cw[251] ^ cw[253] ^ cw[254] ^ cw[257] ^ cw[259] ^ cw[260] ^ cw[263] ^ cw[265] ^ cw[266] ^ cw[268] ^ cw[271] ^ cw[273] ^ cw[275] ^ cw[277] ^ cw[279] ^ cw[280] ^ cw[283] ^ cw[285] ^ cw[287] ^ cw[289] ^ cw[291] ^ cw[292] ^ cw[295] ^ cw[297] ^ cw[299] ^ cw[301] ^ cw[302] ^ cw[305] ^ cw[307] ^ cw[309] ^ cw[310] ^ cw[313] ^ cw[315] ^ cw[316] ^ cw[319] ^ cw[321] ^ cw[322] ^ cw[324] ^ cw[327] ^ cw[329] ^ cw[331] ^ cw[333] ^ cw[334] ^ cw[337] ^ cw[339] ^ cw[341] ^ cw[343] ^ cw[344] ^ cw[347] ^ cw[349] ^ cw[351] ^ cw[352] ^ cw[355] ^ cw[357] ^ cw[358] ^ cw[361] ^ cw[363] ^ cw[364] ^ cw[366] ^ cw[369] ^ cw[371] ^ cw[373] ^ cw[374] ^ cw[377] ^ cw[379] ^ cw[381] ^ cw[382] ^ cw[385] ^ cw[387] ^ cw[388] ^ cw[391] ^ cw[393] ^ cw[394] ^ cw[396] ^ cw[399] ^ cw[401] ^ cw[402] ^ cw[405] ^ cw[407] ^ cw[408] ^ cw[411] ^ cw[413] ^ cw[414] ^ cw[416] ^ cw[419] ^ cw[420] ^ cw[423] ^ cw[425] ^ cw[426] ^ cw[428] ^ cw[431] ^ cw[432] ^ cw[434] ^ cw[437] ^ cw[438] ^ cw[441] ^ cw[443] ^ cw[445] ^ cw[447] ^ cw[449] ^ cw[450] ^ cw[453] ^ cw[455] ^ cw[457] ^ cw[459] ^ cw[461] ^ cw[463] ^ cw[464] ^ cw[467] ^ cw[469] ^ cw[471] ^ cw[473] ^ cw[475] ^ cw[476] ^ cw[479] ^ cw[481] ^ cw[483] ^ cw[485] ^ cw[486] ^ cw[489] ^ cw[491] ^ cw[493] ^ cw[494] ^ cw[497] ^ cw[499] ^ cw[500] ^ cw[503] ^ cw[505] ^ cw[506] ^ cw[508] ^ cw[511] ^ cw[513] ^ cw[515] ^ cw[517] ^ cw[519] ^ cw[520] ^ cw[523] ^ cw[525] ^ cw[527] ^ cw[529] ^ cw[531] ^ cw[532] ^ cw[535] ^ cw[537] ^ cw[539] ^ cw[541] ^ cw[542] ^ cw[545] ^ cw[547] ^ cw[549] ^ cw[550] ^ cw[553] ^ cw[555] ^ cw[556] ^ cw[559] ^ cw[561] ^ cw[562] ^ cw[564] ^ cw[567] ^ cw[569] ^ cw[571] ^ cw[573] ^ cw[574] ^ cw[577] ^ cw[579] ^ cw[581] ^ cw[583] ^ cw[584] ^ cw[587] ^ cw[589] ^ cw[591] ^ cw[592] ^ cw[595] ^ cw[597] ^ cw[598] ^ cw[601] ^ cw[603] ^ cw[604] ^ cw[606] ^ cw[609] ^ cw[611] ^ cw[613] ^ cw[614] ^ cw[617] ^ cw[619] ^ cw[621] ^ cw[622] ^ cw[625] ^ cw[627] ^ cw[628] ^ cw[631] ^ cw[633] ^ cw[634] ^ cw[636] ^ cw[639] ^ cw[641] ^ cw[642] ^ cw[645] ^ cw[647] ^ cw[648] ^ cw[651] ^ cw[653] ^ cw[654] ^ cw[656] ^ cw[659] ^ cw[660] ^ cw[663] ^ cw[665] ^ cw[666] ^ cw[668] ^ cw[671] ^ cw[672] ^ cw[674] ^ cw[677] ^ cw[678] ^ cw[681] ^ cw[683] ^ cw[685] ^ cw[687] ^ cw[688] ^ cw[691] ^ cw[693] ^ cw[695] ^ cw[697] ^ cw[699] ^ cw[700] ^ cw[703] ^ cw[705] ^ cw[707] ^ cw[709] ^ cw[710] ^ cw[713] ^ cw[715] ^ cw[717] ^ cw[718] ^ cw[721] ^ cw[723] ^ cw[724] ^ cw[727] ^ cw[729] ^ cw[730] ^ cw[732] ^ cw[735] ^ cw[737] ^ cw[739] ^ cw[741] ^ cw[742] ^ cw[745] ^ cw[747] ^ cw[749] ^ cw[751] ^ cw[752] ^ cw[755] ^ cw[757] ^ cw[759] ^ cw[760] ^ cw[763] ^ cw[765] ^ cw[766] ^ cw[769] ^ cw[771] ^ cw[772] ^ cw[774] ^ cw[777] ^ cw[779] ^ cw[781] ^ cw[782] ^ cw[785] ^ cw[787] ^ cw[789] ^ cw[790] ^ cw[793] ^ cw[795] ^ cw[796] ^ cw[799] ^ cw[801] ^ cw[802] ^ cw[804] ^ cw[807] ^ cw[809] ^ cw[810] ^ cw[813] ^ cw[815] ^ cw[816] ^ cw[819] ^ cw[821] ^ cw[822] ^ cw[824] ^ cw[827] ^ cw[828] ^ cw[831] ^ cw[833] ^ cw[834] ^ cw[836] ^ cw[839] ^ cw[840] ^ cw[842] ^ cw[845] ^ cw[846] ^ cw[849] ^ cw[851] ^ cw[853] ^ cw[854] ^ cw[857] ^ cw[859] ^ cw[861] ^ cw[863] ^ cw[864] ^ cw[867] ^ cw[869] ^ cw[871] ^ cw[872] ^ cw[875] ^ cw[877] ^ cw[878] ^ cw[881] ^ cw[883] ^ cw[884] ^ cw[886] ^ cw[889] ^ cw[891] ^ cw[893] ^ cw[894] ^ cw[897] ^ cw[899] ^ cw[901] ^ cw[902] ^ cw[905] ^ cw[907] ^ cw[908] ^ cw[911] ^ cw[913] ^ cw[914] ^ cw[916] ^ cw[919] ^ cw[921] ^ cw[922] ^ cw[925] ^ cw[927] ^ cw[928] ^ cw[931] ^ cw[933] ^ cw[934] ^ cw[936] ^ cw[939] ^ cw[940] ^ cw[943] ^ cw[945] ^ cw[946] ^ cw[948] ^ cw[951] ^ cw[952] ^ cw[954] ^ cw[957] ^ cw[958] ^ cw[961] ^ cw[963] ^ cw[964] ^ cw[967] ^ cw[969] ^ cw[971] ^ cw[972] ^ cw[975] ^ cw[977] ^ cw[978] ^ cw[981] ^ cw[983] ^ cw[984] ^ cw[986] ^ cw[989] ^ cw[991] ^ cw[992] ^ cw[995] ^ cw[997] ^ cw[998] ^ cw[1001] ^ cw[1003] ^ cw[1004] ^ cw[1006] ^ cw[1009] ^ cw[1010] ^ cw[1013] ^ cw[1015] ^ cw[1016] ^ cw[1018] ^ cw[1021] ^ cw[1022] ^ cw[1024] ^ cw[1027] ^ cw[1028] ^ cw[1031] ^ cw[1032] ^ cw[1035] ^ cw[1037] ^ cw[1038] ^ cw[1041] ^ cw[1043] ^ cw[1044] ^ cw[1046] ^ cw[1049] ^ cw[1050] ^ cw[1053] ^ cw[1055] ^ cw[1056] ^ cw[1058] ^ cw[1061] ^ cw[1062] ^ cw[1064] ^ cw[1067] ^ cw[1068] ^ cw[1070] ^ cw[1073] ^ cw[1075] ^ cw[1076] ^ cw[1078] ^ cw[1081] ^ cw[1082] ^ cw[1084] ^ cw[1087] ^ cw[1088] ^ cw[1090] ^ cw[1092] ^ cw[1095] ^ cw[1096] ^ cw[1098] ^ cw[1101] ^ cw[1103] ^ cw[1105] ^ cw[1107] ^ cw[1108] ^ cw[1111] ^ cw[1113] ^ cw[1115] ^ cw[1117] ^ cw[1119] ^ cw[1120] ^ cw[1123] ^ cw[1125] ^ cw[1127] ^ cw[1129] ^ cw[1130] ^ cw[1133] ^ cw[1135] ^ cw[1137] ^ cw[1138] ^ cw[1141] ^ cw[1143] ^ cw[1144] ^ cw[1147] ^ cw[1149] ^ cw[1150] ^ cw[1152] ^ cw[1155] ^ cw[1157] ^ cw[1159] ^ cw[1161] ^ cw[1162] ^ cw[1165] ^ cw[1167] ^ cw[1169] ^ cw[1171] ^ cw[1172] ^ cw[1175] ^ cw[1177] ^ cw[1179] ^ cw[1180] ^ cw[1183] ^ cw[1185] ^ cw[1186] ^ cw[1189] ^ cw[1191] ^ cw[1192] ^ cw[1194] ^ cw[1197] ^ cw[1199] ^ cw[1201] ^ cw[1202] ^ cw[1205] ^ cw[1207] ^ cw[1209] ^ cw[1210] ^ cw[1213] ^ cw[1215] ^ cw[1216] ^ cw[1219] ^ cw[1221] ^ cw[1222] ^ cw[1224] ^ cw[1227] ^ cw[1229] ^ cw[1230] ^ cw[1233] ^ cw[1235] ^ cw[1236] ^ cw[1239] ^ cw[1241] ^ cw[1242] ^ cw[1244] ^ cw[1247] ^ cw[1248] ^ cw[1251] ^ cw[1253] ^ cw[1254] ^ cw[1256] ^ cw[1259] ^ cw[1260] ^ cw[1262] ^ cw[1265] ^ cw[1266] ^ cw[1269] ^ cw[1271] ^ cw[1273] ^ cw[1274] ^ cw[1277] ^ cw[1279] ^ cw[1281] ^ cw[1283] ^ cw[1284] ^ cw[1287] ^ cw[1289] ^ cw[1291] ^ cw[1292] ^ cw[1295] ^ cw[1297] ^ cw[1298] ^ cw[1301] ^ cw[1303] ^ cw[1304] ^ cw[1306] ^ cw[1309] ^ cw[1311] ^ cw[1313] ^ cw[1314] ^ cw[1317] ^ cw[1319] ^ cw[1321] ^ cw[1322] ^ cw[1325] ^ cw[1327] ^ cw[1328] ^ cw[1331] ^ cw[1333] ^ cw[1334] ^ cw[1336] ^ cw[1339] ^ cw[1341] ^ cw[1342] ^ cw[1345] ^ cw[1347] ^ cw[1348] ^ cw[1351] ^ cw[1353] ^ cw[1354] ^ cw[1356] ^ cw[1359] ^ cw[1360] ^ cw[1363] ^ cw[1365] ^ cw[1366] ^ cw[1368] ^ cw[1371] ^ cw[1372] ^ cw[1374] ^ cw[1377] ^ cw[1378] ^ cw[1381] ^ cw[1383] ^ cw[1384] ^ cw[1387] ^ cw[1389] ^ cw[1391] ^ cw[1392] ^ cw[1395] ^ cw[1397] ^ cw[1398] ^ cw[1401] ^ cw[1403] ^ cw[1404] ^ cw[1406] ^ cw[1409] ^ cw[1411] ^ cw[1412] ^ cw[1415] ^ cw[1417] ^ cw[1418] ^ cw[1421] ^ cw[1423] ^ cw[1424] ^ cw[1426] ^ cw[1429] ^ cw[1430] ^ cw[1433] ^ cw[1435] ^ cw[1436] ^ cw[1438] ^ cw[1441] ^ cw[1442] ^ cw[1444] ^ cw[1447] ^ cw[1448] ^ cw[1451] ^ cw[1452] ^ cw[1455] ^ cw[1457] ^ cw[1458] ^ cw[1461] ^ cw[1463] ^ cw[1464] ^ cw[1466] ^ cw[1469] ^ cw[1470] ^ cw[1473] ^ cw[1475] ^ cw[1476] ^ cw[1478] ^ cw[1481] ^ cw[1482] ^ cw[1484] ^ cw[1487] ^ cw[1488] ^ cw[1490] ^ cw[1493] ^ cw[1495] ^ cw[1496] ^ cw[1498] ^ cw[1501] ^ cw[1502] ^ cw[1504] ^ cw[1507] ^ cw[1508] ^ cw[1510] ^ cw[1512] ^ cw[1515] ^ cw[1516] ^ cw[1518] ^ cw[1521] ^ cw[1523] ^ cw[1525] ^ cw[1526] ^ cw[1529] ^ cw[1531] ^ cw[1533] ^ cw[1535] ^ cw[1536] ^ cw[1539] ^ cw[1541] ^ cw[1543] ^ cw[1544] ^ cw[1547] ^ cw[1549] ^ cw[1550] ^ cw[1553] ^ cw[1555] ^ cw[1556] ^ cw[1558] ^ cw[1561] ^ cw[1563] ^ cw[1565] ^ cw[1566] ^ cw[1569] ^ cw[1571] ^ cw[1573] ^ cw[1574] ^ cw[1577] ^ cw[1579] ^ cw[1580] ^ cw[1583] ^ cw[1585] ^ cw[1586] ^ cw[1588] ^ cw[1591] ^ cw[1593] ^ cw[1594] ^ cw[1597] ^ cw[1599] ^ cw[1600] ^ cw[1603] ^ cw[1605] ^ cw[1606] ^ cw[1608] ^ cw[1611] ^ cw[1612] ^ cw[1615] ^ cw[1617] ^ cw[1618] ^ cw[1620] ^ cw[1623] ^ cw[1624] ^ cw[1626] ^ cw[1629] ^ cw[1630] ^ cw[1633] ^ cw[1635] ^ cw[1636] ^ cw[1639] ^ cw[1641] ^ cw[1643] ^ cw[1644] ^ cw[1647] ^ cw[1649] ^ cw[1650] ^ cw[1653] ^ cw[1655] ^ cw[1656] ^ cw[1658] ^ cw[1661] ^ cw[1663] ^ cw[1664] ^ cw[1667] ^ cw[1669] ^ cw[1670] ^ cw[1673] ^ cw[1675] ^ cw[1676] ^ cw[1678] ^ cw[1681] ^ cw[1682] ^ cw[1685] ^ cw[1687] ^ cw[1688] ^ cw[1690] ^ cw[1693] ^ cw[1694] ^ cw[1696] ^ cw[1699] ^ cw[1700] ^ cw[1703] ^ cw[1704] ^ cw[1707] ^ cw[1709] ^ cw[1710] ^ cw[1713] ^ cw[1715] ^ cw[1716] ^ cw[1718] ^ cw[1721] ^ cw[1722] ^ cw[1725] ^ cw[1727] ^ cw[1728] ^ cw[1730] ^ cw[1733] ^ cw[1734] ^ cw[1736] ^ cw[1739] ^ cw[1740] ^ cw[1742] ^ cw[1745] ^ cw[1747] ^ cw[1748] ^ cw[1750] ^ cw[1753] ^ cw[1754] ^ cw[1756] ^ cw[1759] ^ cw[1760] ^ cw[1762] ^ cw[1764] ^ cw[1767] ^ cw[1768] ^ cw[1770] ^ cw[1773] ^ cw[1775] ^ cw[1776] ^ cw[1779] ^ cw[1781] ^ cw[1783] ^ cw[1784] ^ cw[1787] ^ cw[1789] ^ cw[1790] ^ cw[1793] ^ cw[1795] ^ cw[1796] ^ cw[1798] ^ cw[1801] ^ cw[1803] ^ cw[1804] ^ cw[1807] ^ cw[1809] ^ cw[1810] ^ cw[1813] ^ cw[1815] ^ cw[1816] ^ cw[1818] ^ cw[1821] ^ cw[1822] ^ cw[1825] ^ cw[1827] ^ cw[1828] ^ cw[1830] ^ cw[1833] ^ cw[1834] ^ cw[1836] ^ cw[1839] ^ cw[1840] ^ cw[1843] ^ cw[1844] ^ cw[1847] ^ cw[1849] ^ cw[1850] ^ cw[1853] ^ cw[1855] ^ cw[1856] ^ cw[1858] ^ cw[1861] ^ cw[1862] ^ cw[1865] ^ cw[1867] ^ cw[1868] ^ cw[1870] ^ cw[1873] ^ cw[1874] ^ cw[1876] ^ cw[1879] ^ cw[1880] ^ cw[1882] ^ cw[1885] ^ cw[1887] ^ cw[1888] ^ cw[1890] ^ cw[1893] ^ cw[1894] ^ cw[1896] ^ cw[1899] ^ cw[1900] ^ cw[1902] ^ cw[1904] ^ cw[1907] ^ cw[1908] ^ cw[1910] ^ cw[1913] ^ cw[1914] ^ cw[1917] ^ cw[1919] ^ cw[1920] ^ cw[1923] ^ cw[1925] ^ cw[1926] ^ cw[1928] ^ cw[1931] ^ cw[1932] ^ cw[1935] ^ cw[1937] ^ cw[1938] ^ cw[1940] ^ cw[1943] ^ cw[1944] ^ cw[1946] ^ cw[1949] ^ cw[1950] ^ cw[1952] ^ cw[1955] ^ cw[1957] ^ cw[1958] ^ cw[1960] ^ cw[1963] ^ cw[1964] ^ cw[1966] ^ cw[1969] ^ cw[1970] ^ cw[1972] ^ cw[1974] ^ cw[1977] ^ cw[1978] ^ cw[1980] ^ cw[1982] ^ cw[1985] ^ cw[1987] ^ cw[1988] ^ cw[1990] ^ cw[1993] ^ cw[1994] ^ cw[1996] ^ cw[1999] ^ cw[2000] ^ cw[2002] ^ cw[2004] ^ cw[2007] ^ cw[2008] ^ cw[2010] ^ cw[2012] ^ cw[2014] ^ cw[2017] ^ cw[2018] ^ cw[2020] ^ cw[2022] ^ cw[2024] ^ cw[2025] ^ cw[2027] ^ cw[2028] ^ cw[2029] ^ cw[2030] ^ cw[2031] ^ cw[2032] ^ cw[2033] ^ cw[2034] ^ cw[2035] ^ cw[2038];
    assign syndrome[8] = cw[1] ^ cw[3] ^ cw[5] ^ cw[7] ^ cw[9] ^ cw[11] ^ cw[12] ^ cw[15] ^ cw[17] ^ cw[19] ^ cw[21] ^ cw[23] ^ cw[25] ^ cw[27] ^ cw[29] ^ cw[30] ^ cw[33] ^ cw[35] ^ cw[37] ^ cw[39] ^ cw[41] ^ cw[43] ^ cw[45] ^ cw[46] ^ cw[49] ^ cw[51] ^ cw[53] ^ cw[55] ^ cw[57] ^ cw[59] ^ cw[60] ^ cw[63] ^ cw[65] ^ cw[67] ^ cw[69] ^ cw[71] ^ cw[72] ^ cw[75] ^ cw[77] ^ cw[79] ^ cw[81] ^ cw[82] ^ cw[85] ^ cw[87] ^ cw[89] ^ cw[90] ^ cw[93] ^ cw[95] ^ cw[97] ^ cw[98] ^ cw[100] ^ cw[102] ^ cw[105] ^ cw[107] ^ cw[109] ^ cw[111] ^ cw[113] ^ cw[115] ^ cw[117] ^ cw[119] ^ cw[120] ^ cw[123] ^ cw[125] ^ cw[127] ^ cw[129] ^ cw[131] ^ cw[133] ^ cw[135] ^ cw[136] ^ cw[139] ^ cw[141] ^ cw[143] ^ cw[145] ^ cw[147] ^ cw[149] ^ cw[150] ^ cw[153] ^ cw[155] ^ cw[157] ^ cw[159] ^ cw[161] ^ cw[162] ^ cw[165] ^ cw[167] ^ cw[169] ^ cw[171] ^ cw[172] ^ cw[175] ^ cw[177] ^ cw[179] ^ cw[180] ^ cw[183] ^ cw[185] ^ cw[187] ^ cw[188] ^ cw[190] ^ cw[192] ^ cw[195] ^ cw[197] ^ cw[199] ^ cw[201] ^ cw[203] ^ cw[205] ^ cw[207] ^ cw[208] ^ cw[211] ^ cw[213] ^ cw[215] ^ cw[217] ^ cw[219] ^ cw[221] ^ cw[222] ^ cw[225] ^ cw[227] ^ cw[229] ^ cw[231] ^ cw[233] ^ cw[234] ^ cw[237] ^ cw[239] ^ cw[241] ^ cw[243] ^ cw[244] ^ cw[247] ^ cw[249] ^ cw[251] ^ cw[252] ^ cw[255] ^ cw[257] ^ cw[259] ^ cw[260] ^ cw[262] ^ cw[264] ^ cw[267] ^ cw[269] ^ cw[271] ^ cw[273] ^ cw[275] ^ cw[277] ^ cw[278] ^ cw[281] ^ cw[283] ^ cw[285] ^ cw[287] ^ cw[289] ^ cw[290] ^ cw[293] ^ cw[295] ^ cw[297] ^ cw[299] ^ cw[300] ^ cw[303] ^ cw[305] ^ cw[307] ^ cw[308] ^ cw[311] ^ cw[313] ^ cw[315] ^ cw[316] ^ cw[318] ^ cw[320] ^ cw[323] ^ cw[325] ^ cw[327] ^ cw[329] ^ cw[331] ^ cw[332] ^ cw[335] ^ cw[337] ^ cw[339] ^ cw[341] ^ cw[342] ^ cw[345] ^ cw[347] ^ cw[349] ^ cw[350] ^ cw[353] ^ cw[355] ^ cw[357] ^ cw[358] ^ cw[360] ^ cw[362] ^ cw[365] ^ cw[367] ^ cw[369] ^ cw[371] ^ cw[372] ^ cw[375] ^ cw[377] ^ cw[379] ^ cw[380] ^ cw[383] ^ cw[385] ^ cw[387] ^ cw[388] ^ cw[390] ^ cw[392] ^ cw[395] ^ cw[397] ^ cw[399] ^ cw[400] ^ cw[403] ^ cw[405] ^ cw[407] ^ cw[408] ^ cw[410] ^ cw[412] ^ cw[415] ^ cw[417] ^ cw[419] ^ cw[420] ^ cw[422] ^ cw[424] ^ cw[427] ^ cw[429] ^ cw[431] ^ cw[432] ^ cw[434] ^ cw[436] ^ cw[439] ^ cw[441] ^ cw[443] ^ cw[445] ^ cw[447] ^ cw[448] ^ cw[451] ^ cw[453] ^ cw[455] ^ cw[457] ^ cw[459] ^ cw[461] ^ cw[462] ^ cw[465] ^ cw[467] ^ cw[469] ^ cw[471] ^ cw[473] ^ cw[474] ^ cw[477] ^ cw[479] ^ cw[481] ^ cw[483] ^ cw[484] ^ cw[487] ^ cw[489] ^ cw[491] ^ cw[492] ^ cw[495] ^ cw[497] ^ cw[499] ^ cw[500] ^ cw[502] ^ cw[504] ^ cw[507] ^ cw[509] ^ cw[511] ^ cw[513] ^ cw[515] ^ cw[517] ^ cw[518] ^ cw[521] ^ cw[523] ^ cw[525] ^ cw[527] ^ cw[529] ^ cw[530] ^ cw[533] ^ cw[535] ^ cw[537] ^ cw[539] ^ cw[540] ^ cw[543] ^ cw[545] ^ cw[547] ^ cw[548] ^ cw[551] ^ cw[553] ^ cw[555] ^ cw[556] ^ cw[558] ^ cw[560] ^ cw[563] ^ cw[565] ^ cw[567] ^ cw[569] ^ cw[571] ^ cw[572] ^ cw[575] ^ cw[577] ^ cw[579] ^ cw[581] ^ cw[582] ^ cw[585] ^ cw[587] ^ cw[589] ^ cw[590] ^ cw[593] ^ cw[595] ^ cw[597] ^ cw[598] ^ cw[600] ^ cw[602] ^ cw[605] ^ cw[607] ^ cw[609] ^ cw[611] ^ cw[612] ^ cw[615] ^ cw[617] ^ cw[619] ^ cw[620] ^ cw[623] ^ cw[625] ^ cw[627] ^ cw[628] ^ cw[630] ^ cw[632] ^ cw[635] ^ cw[637] ^ cw[639] ^ cw[640] ^ cw[643] ^ cw[645] ^ cw[647] ^ cw[648] ^ cw[650] ^ cw[652] ^ cw[655] ^ cw[657] ^ cw[659] ^ cw[660] ^ cw[662] ^ cw[664] ^ cw[667] ^ cw[669] ^ cw[671] ^ cw[672] ^ cw[674] ^ cw[676] ^ cw[679] ^ cw[681] ^ cw[683] ^ cw[685] ^ cw[686] ^ cw[689] ^ cw[691] ^ cw[693] ^ cw[695] ^ cw[697] ^ cw[698] ^ cw[701] ^ cw[703] ^ cw[705] ^ cw[707] ^ cw[708] ^ cw[711] ^ cw[713] ^ cw[715] ^ cw[716] ^ cw[719] ^ cw[721] ^ cw[723] ^ cw[724] ^ cw[726] ^ cw[728] ^ cw[731] ^ cw[733] ^ cw[735] ^ cw[737] ^ cw[739] ^ cw[740] ^ cw[743] ^ cw[745] ^ cw[747] ^ cw[749] ^ cw[750] ^ cw[753] ^ cw[755] ^ cw[757] ^ cw[758] ^ cw[761] ^ cw[763] ^ cw[765] ^ cw[766] ^ cw[768] ^ cw[770] ^ cw[773] ^ cw[775] ^ cw[777] ^ cw[779] ^ cw[780] ^ cw[783] ^ cw[785] ^ cw[787] ^ cw[788] ^ cw[791] ^ cw[793] ^ cw[795] ^ cw[796] ^ cw[798] ^ cw[800] ^ cw[803] ^ cw[805] ^ cw[807] ^ cw[808] ^ cw[811] ^ cw[813] ^ cw[815] ^ cw[816] ^ cw[818] ^ cw[820] ^ cw[823] ^ cw[825] ^ cw[827] ^ cw[828] ^ cw[830] ^ cw[832] ^ cw[835] ^ cw[837] ^ cw[839] ^ cw[840] ^ cw[842] ^ cw[844] ^ cw[847] ^ cw[849] ^ cw[851] ^ cw[852] ^ cw[855] ^ cw[857] ^ cw[859] ^ cw[861] ^ cw[862] ^ cw[865] ^ cw[867] ^ cw[869] ^ cw[870] ^ cw[873] ^ cw[875] ^ cw[877] ^ cw[878] ^ cw[880] ^ cw[882] ^ cw[885] ^ cw[887] ^ cw[889] ^ cw[891] ^ cw[892] ^ cw[895] ^ cw[897] ^ cw[899] ^ cw[900] ^ cw[903] ^ cw[905] ^ cw[907] ^ cw[908] ^ cw[910] ^ cw[912] ^ cw[915] ^ cw[917] ^ cw[919] ^ cw[920] ^ cw[923] ^ cw[925] ^ cw[927] ^ cw[928] ^ cw[930] ^ cw[932] ^ cw[935] ^ cw[937] ^ cw[939] ^ cw[940] ^ cw[942] ^ cw[944] ^ cw[947] ^ cw[949] ^ cw[951] ^ cw[952] ^ cw[954] ^ cw[956] ^ cw[959] ^ cw[961] ^ cw[962] ^ cw[965] ^ cw[967] ^ cw[969] ^ cw[970] ^ cw[973] ^ cw[975] ^ cw[977] ^ cw[978] ^ cw[980] ^ cw[982] ^ cw[985] ^ cw[987] ^ cw[989] ^ cw[990] ^ cw[993] ^ cw[995] ^ cw[997] ^ cw[998] ^ cw[1000] ^ cw[1002] ^ cw[1005] ^ cw[1007] ^ cw[1009] ^ cw[1010] ^ cw[1012] ^ cw[1014] ^ cw[1017] ^ cw[1019] ^ cw[1021] ^ cw[1022] ^ cw[1024] ^ cw[1026] ^ cw[1029] ^ cw[1030] ^ cw[1033] ^ cw[1035] ^ cw[1037] ^ cw[1038] ^ cw[1040] ^ cw[1042] ^ cw[1045] ^ cw[1047] ^ cw[1049] ^ cw[1050] ^ cw[1052] ^ cw[1054] ^ cw[1057] ^ cw[1059] ^ cw[1061] ^ cw[1062] ^ cw[1064] ^ cw[1066] ^ cw[1069] ^ cw[1070] ^ cw[1072] ^ cw[1074] ^ cw[1077] ^ cw[1079] ^ cw[1081] ^ cw[1082] ^ cw[1084] ^ cw[1086] ^ cw[1089] ^ cw[1090] ^ cw[1092] ^ cw[1094] ^ cw[1097] ^ cw[1098] ^ cw[1101] ^ cw[1103] ^ cw[1105] ^ cw[1106] ^ cw[1109] ^ cw[1111] ^ cw[1113] ^ cw[1115] ^ cw[1117] ^ cw[1118] ^ cw[1121] ^ cw[1123] ^ cw[1125] ^ cw[1127] ^ cw[1128] ^ cw[1131] ^ cw[1133] ^ cw[1135] ^ cw[1136] ^ cw[1139] ^ cw[1141] ^ cw[1143] ^ cw[1144] ^ cw[1146] ^ cw[1148] ^ cw[1151] ^ cw[1153] ^ cw[1155] ^ cw[1157] ^ cw[1159] ^ cw[1160] ^ cw[1163] ^ cw[1165] ^ cw[1167] ^ cw[1169] ^ cw[1170] ^ cw[1173] ^ cw[1175] ^ cw[1177] ^ cw[1178] ^ cw[1181] ^ cw[1183] ^ cw[1185] ^ cw[1186] ^ cw[1188] ^ cw[1190] ^ cw[1193] ^ cw[1195] ^ cw[1197] ^ cw[1199] ^ cw[1200] ^ cw[1203] ^ cw[1205] ^ cw[1207] ^ cw[1208] ^ cw[1211] ^ cw[1213] ^ cw[1215] ^ cw[1216] ^ cw[1218] ^ cw[1220] ^ cw[1223] ^ cw[1225] ^ cw[1227] ^ cw[1228] ^ cw[1231] ^ cw[1233] ^ cw[1235] ^ cw[1236] ^ cw[1238] ^ cw[1240] ^ cw[1243] ^ cw[1245] ^ cw[1247] ^ cw[1248] ^ cw[1250] ^ cw[1252] ^ cw[1255] ^ cw[1257] ^ cw[1259] ^ cw[1260] ^ cw[1262] ^ cw[1264] ^ cw[1267] ^ cw[1269] ^ cw[1271] ^ cw[1272] ^ cw[1275] ^ cw[1277] ^ cw[1279] ^ cw[1281] ^ cw[1282] ^ cw[1285] ^ cw[1287] ^ cw[1289] ^ cw[1290] ^ cw[1293] ^ cw[1295] ^ cw[1297] ^ cw[1298] ^ cw[1300] ^ cw[1302] ^ cw[1305] ^ cw[1307] ^ cw[1309] ^ cw[1311] ^ cw[1312] ^ cw[1315] ^ cw[1317] ^ cw[1319] ^ cw[1320] ^ cw[1323] ^ cw[1325] ^ cw[1327] ^ cw[1328] ^ cw[1330] ^ cw[1332] ^ cw[1335] ^ cw[1337] ^ cw[1339] ^ cw[1340] ^ cw[1343] ^ cw[1345] ^ cw[1347] ^ cw[1348] ^ cw[1350] ^ cw[1352] ^ cw[1355] ^ cw[1357] ^ cw[1359] ^ cw[1360] ^ cw[1362] ^ cw[1364] ^ cw[1367] ^ cw[1369] ^ cw[1371] ^ cw[1372] ^ cw[1374] ^ cw[1376] ^ cw[1379] ^ cw[1381] ^ cw[1382] ^ cw[1385] ^ cw[1387] ^ cw[1389] ^ cw[1390] ^ cw[1393] ^ cw[1395] ^ cw[1397] ^ cw[1398] ^ cw[1400] ^ cw[1402] ^ cw[1405] ^ cw[1407] ^ cw[1409] ^ cw[1410] ^ cw[1413] ^ cw[1415] ^ cw[1417] ^ cw[1418] ^ cw[1420] ^ cw[1422] ^ cw[1425] ^ cw[1427] ^ cw[1429] ^ cw[1430] ^ cw[1432] ^ cw[1434] ^ cw[1437] ^ cw[1439] ^ cw[1441] ^ cw[1442] ^ cw[1444] ^ cw[1446] ^ cw[1449] ^ cw[1450] ^ cw[1453] ^ cw[1455] ^ cw[1457] ^ cw[1458] ^ cw[1460] ^ cw[1462] ^ cw[1465] ^ cw[1467] ^ cw[1469] ^ cw[1470] ^ cw[1472] ^ cw[1474] ^ cw[1477] ^ cw[1479] ^ cw[1481] ^ cw[1482] ^ cw[1484] ^ cw[1486] ^ cw[1489] ^ cw[1490] ^ cw[1492] ^ cw[1494] ^ cw[1497] ^ cw[1499] ^ cw[1501] ^ cw[1502] ^ cw[1504] ^ cw[1506] ^ cw[1509] ^ cw[1510] ^ cw[1512] ^ cw[1514] ^ cw[1517] ^ cw[1518] ^ cw[1521] ^ cw[1523] ^ cw[1524] ^ cw[1527] ^ cw[1529] ^ cw[1531] ^ cw[1533] ^ cw[1534] ^ cw[1537] ^ cw[1539] ^ cw[1541] ^ cw[1542] ^ cw[1545] ^ cw[1547] ^ cw[1549] ^ cw[1550] ^ cw[1552] ^ cw[1554] ^ cw[1557] ^ cw[1559] ^ cw[1561] ^ cw[1563] ^ cw[1564] ^ cw[1567] ^ cw[1569] ^ cw[1571] ^ cw[1572] ^ cw[1575] ^ cw[1577] ^ cw[1579] ^ cw[1580] ^ cw[1582] ^ cw[1584] ^ cw[1587] ^ cw[1589] ^ cw[1591] ^ cw[1592] ^ cw[1595] ^ cw[1597] ^ cw[1599] ^ cw[1600] ^ cw[1602] ^ cw[1604] ^ cw[1607] ^ cw[1609] ^ cw[1611] ^ cw[1612] ^ cw[1614] ^ cw[1616] ^ cw[1619] ^ cw[1621] ^ cw[1623] ^ cw[1624] ^ cw[1626] ^ cw[1628] ^ cw[1631] ^ cw[1633] ^ cw[1634] ^ cw[1637] ^ cw[1639] ^ cw[1641] ^ cw[1642] ^ cw[1645] ^ cw[1647] ^ cw[1649] ^ cw[1650] ^ cw[1652] ^ cw[1654] ^ cw[1657] ^ cw[1659] ^ cw[1661] ^ cw[1662] ^ cw[1665] ^ cw[1667] ^ cw[1669] ^ cw[1670] ^ cw[1672] ^ cw[1674] ^ cw[1677] ^ cw[1679] ^ cw[1681] ^ cw[1682] ^ cw[1684] ^ cw[1686] ^ cw[1689] ^ cw[1691] ^ cw[1693] ^ cw[1694] ^ cw[1696] ^ cw[1698] ^ cw[1701] ^ cw[1702] ^ cw[1705] ^ cw[1707] ^ cw[1709] ^ cw[1710] ^ cw[1712] ^ cw[1714] ^ cw[1717] ^ cw[1719] ^ cw[1721] ^ cw[1722] ^ cw[1724] ^ cw[1726] ^ cw[1729] ^ cw[1731] ^ cw[1733] ^ cw[1734] ^ cw[1736] ^ cw[1738] ^ cw[1741] ^ cw[1742] ^ cw[1744] ^ cw[1746] ^ cw[1749] ^ cw[1751] ^ cw[1753] ^ cw[1754] ^ cw[1756] ^ cw[1758] ^ cw[1761] ^ cw[1762] ^ cw[1764] ^ cw[1766] ^ cw[1769] ^ cw[1770] ^ cw[1773] ^ cw[1774] ^ cw[1777] ^ cw[1779] ^ cw[1781] ^ cw[1782] ^ cw[1785] ^ cw[1787] ^ cw[1789] ^ cw[1790] ^ cw[1792] ^ cw[1794] ^ cw[1797] ^ cw[1799] ^ cw[1801] ^ cw[1802] ^ cw[1805] ^ cw[1807] ^ cw[1809] ^ cw[1810] ^ cw[1812] ^ cw[1814] ^ cw[1817] ^ cw[1819] ^ cw[1821] ^ cw[1822] ^ cw[1824] ^ cw[1826] ^ cw[1829] ^ cw[1831] ^ cw[1833] ^ cw[1834] ^ cw[1836] ^ cw[1838] ^ cw[1841] ^ cw[1842] ^ cw[1845] ^ cw[1847] ^ cw[1849] ^ cw[1850] ^ cw[1852] ^ cw[1854] ^ cw[1857] ^ cw[1859] ^ cw[1861] ^ cw[1862] ^ cw[1864] ^ cw[1866] ^ cw[1869] ^ cw[1871] ^ cw[1873] ^ cw[1874] ^ cw[1876] ^ cw[1878] ^ cw[1881] ^ cw[1882] ^ cw[1884] ^ cw[1886] ^ cw[1889] ^ cw[1891] ^ cw[1893] ^ cw[1894] ^ cw[1896] ^ cw[1898] ^ cw[1901] ^ cw[1902] ^ cw[1904] ^ cw[1906] ^ cw[1909] ^ cw[1910] ^ cw[1912] ^ cw[1915] ^ cw[1917] ^ cw[1919] ^ cw[1920] ^ cw[1922] ^ cw[1924] ^ cw[1927] ^ cw[1929] ^ cw[1931] ^ cw[1932] ^ cw[1934] ^ cw[1936] ^ cw[1939] ^ cw[1941] ^ cw[1943] ^ cw[1944] ^ cw[1946] ^ cw[1948] ^ cw[1951] ^ cw[1952] ^ cw[1954] ^ cw[1956] ^ cw[1959] ^ cw[1961] ^ cw[1963] ^ cw[1964] ^ cw[1966] ^ cw[1968] ^ cw[1971] ^ cw[1972] ^ cw[1974] ^ cw[1976] ^ cw[1979] ^ cw[1980] ^ cw[1982] ^ cw[1984] ^ cw[1986] ^ cw[1989] ^ cw[1991] ^ cw[1993] ^ cw[1994] ^ cw[1996] ^ cw[1998] ^ cw[2001] ^ cw[2002] ^ cw[2004] ^ cw[2006] ^ cw[2009] ^ cw[2010] ^ cw[2012] ^ cw[2014] ^ cw[2016] ^ cw[2019] ^ cw[2020] ^ cw[2022] ^ cw[2024] ^ cw[2025] ^ cw[2026] ^ cw[2028] ^ cw[2029] ^ cw[2030] ^ cw[2031] ^ cw[2032] ^ cw[2033] ^ cw[2034] ^ cw[2035] ^ cw[2039];
    assign syndrome[7] = cw[1] ^ cw[3] ^ cw[5] ^ cw[7] ^ cw[9] ^ cw[10] ^ cw[13] ^ cw[15] ^ cw[17] ^ cw[19] ^ cw[21] ^ cw[23] ^ cw[25] ^ cw[27] ^ cw[28] ^ cw[31] ^ cw[33] ^ cw[35] ^ cw[37] ^ cw[39] ^ cw[41] ^ cw[43] ^ cw[44] ^ cw[47] ^ cw[49] ^ cw[51] ^ cw[53] ^ cw[55] ^ cw[57] ^ cw[58] ^ cw[61] ^ cw[63] ^ cw[65] ^ cw[67] ^ cw[69] ^ cw[70] ^ cw[73] ^ cw[75] ^ cw[77] ^ cw[79] ^ cw[80] ^ cw[83] ^ cw[85] ^ cw[87] ^ cw[89] ^ cw[90] ^ cw[92] ^ cw[94] ^ cw[96] ^ cw[99] ^ cw[101] ^ cw[103] ^ cw[105] ^ cw[107] ^ cw[109] ^ cw[111] ^ cw[113] ^ cw[115] ^ cw[117] ^ cw[118] ^ cw[121] ^ cw[123] ^ cw[125] ^ cw[127] ^ cw[129] ^ cw[131] ^ cw[133] ^ cw[134] ^ cw[137] ^ cw[139] ^ cw[141] ^ cw[143] ^ cw[145] ^ cw[147] ^ cw[148] ^ cw[151] ^ cw[153] ^ cw[155] ^ cw[157] ^ cw[159] ^ cw[160] ^ cw[163] ^ cw[165] ^ cw[167] ^ cw[169] ^ cw[170] ^ cw[173] ^ cw[175] ^ cw[177] ^ cw[179] ^ cw[180] ^ cw[182] ^ cw[184] ^ cw[186] ^ cw[189] ^ cw[191] ^ cw[193] ^ cw[195] ^ cw[197] ^ cw[199] ^ cw[201] ^ cw[203] ^ cw[205] ^ cw[206] ^ cw[209] ^ cw[211] ^ cw[213] ^ cw[215] ^ cw[217] ^ cw[219] ^ cw[220] ^ cw[223] ^ cw[225] ^ cw[227] ^ cw[229] ^ cw[231] ^ cw[232] ^ cw[235] ^ cw[237] ^ cw[239] ^ cw[241] ^ cw[242] ^ cw[245] ^ cw[247] ^ cw[249] ^ cw[251] ^ cw[252] ^ cw[254] ^ cw[256] ^ cw[258] ^ cw[261] ^ cw[263] ^ cw[265] ^ cw[267] ^ cw[269] ^ cw[271] ^ cw[273] ^ cw[275] ^ cw[276] ^ cw[279] ^ cw[281] ^ cw[283] ^ cw[285] ^ cw[287] ^ cw[288] ^ cw[291] ^ cw[293] ^ cw[295] ^ cw[297] ^ cw[298] ^ cw[301] ^ cw[303] ^ cw[305] ^ cw[307] ^ cw[308] ^ cw[310] ^ cw[312] ^ cw[314] ^ cw[317] ^ cw[319] ^ cw[321] ^ cw[323] ^ cw[325] ^ cw[327] ^ cw[329] ^ cw[330] ^ cw[333] ^ cw[335] ^ cw[337] ^ cw[339] ^ cw[340] ^ cw[343] ^ cw[345] ^ cw[347] ^ cw[349] ^ cw[350] ^ cw[352] ^ cw[354] ^ cw[356] ^ cw[359] ^ cw[361] ^ cw[363] ^ cw[365] ^ cw[367] ^ cw[369] ^ cw[370] ^ cw[373] ^ cw[375] ^ cw[377] ^ cw[379] ^ cw[380] ^ cw[382] ^ cw[384] ^ cw[386] ^ cw[389] ^ cw[391] ^ cw[393] ^ cw[395] ^ cw[397] ^ cw[399] ^ cw[400] ^ cw[402] ^ cw[404] ^ cw[406] ^ cw[409] ^ cw[411] ^ cw[413] ^ cw[415] ^ cw[417] ^ cw[419] ^ cw[420] ^ cw[422] ^ cw[424] ^ cw[426] ^ cw[428] ^ cw[430] ^ cw[433] ^ cw[435] ^ cw[437] ^ cw[439] ^ cw[441] ^ cw[443] ^ cw[445] ^ cw[446] ^ cw[449] ^ cw[451] ^ cw[453] ^ cw[455] ^ cw[457] ^ cw[459] ^ cw[460] ^ cw[463] ^ cw[465] ^ cw[467] ^ cw[469] ^ cw[471] ^ cw[472] ^ cw[475] ^ cw[477] ^ cw[479] ^ cw[481] ^ cw[482] ^ cw[485] ^ cw[487] ^ cw[489] ^ cw[491] ^ cw[492] ^ cw[494] ^ cw[496] ^ cw[498] ^ cw[501] ^ cw[503] ^ cw[505] ^ cw[507] ^ cw[509] ^ cw[511] ^ cw[513] ^ cw[515] ^ cw[516] ^ cw[519] ^ cw[521] ^ cw[523] ^ cw[525] ^ cw[527] ^ cw[528] ^ cw[531] ^ cw[533] ^ cw[535] ^ cw[537] ^ cw[538] ^ cw[541] ^ cw[543] ^ cw[545] ^ cw[547] ^ cw[548] ^ cw[550] ^ cw[552] ^ cw[554] ^ cw[557] ^ cw[559] ^ cw[561] ^ cw[563] ^ cw[565] ^ cw[567] ^ cw[569] ^ cw[570] ^ cw[573] ^ cw[575] ^ cw[577] ^ cw[579] ^ cw[580] ^ cw[583] ^ cw[585] ^ cw[587] ^ cw[589] ^ cw[590] ^ cw[592] ^ cw[594] ^ cw[596] ^ cw[599] ^ cw[601] ^ cw[603] ^ cw[605] ^ cw[607] ^ cw[609] ^ cw[610] ^ cw[613] ^ cw[615] ^ cw[617] ^ cw[619] ^ cw[620] ^ cw[622] ^ cw[624] ^ cw[626] ^ cw[629] ^ cw[631] ^ cw[633] ^ cw[635] ^ cw[637] ^ cw[639] ^ cw[640] ^ cw[642] ^ cw[644] ^ cw[646] ^ cw[649] ^ cw[651] ^ cw[653] ^ cw[655] ^ cw[657] ^ cw[659] ^ cw[660] ^ cw[662] ^ cw[664] ^ cw[666] ^ cw[668] ^ cw[670] ^ cw[673] ^ cw[675] ^ cw[677] ^ cw[679] ^ cw[681] ^ cw[683] ^ cw[684] ^ cw[687] ^ cw[689] ^ cw[691] ^ cw[693] ^ cw[695] ^ cw[696] ^ cw[699] ^ cw[701] ^ cw[703] ^ cw[705] ^ cw[706] ^ cw[709] ^ cw[711] ^ cw[713] ^ cw[715] ^ cw[716] ^ cw[718] ^ cw[720] ^ cw[722] ^ cw[725] ^ cw[727] ^ cw[729] ^ cw[731] ^ cw[733] ^ cw[735] ^ cw[737] ^ cw[738] ^ cw[741] ^ cw[743] ^ cw[745] ^ cw[747] ^ cw[748] ^ cw[751] ^ cw[753] ^ cw[755] ^ cw[757] ^ cw[758] ^ cw[760] ^ cw[762] ^ cw[764] ^ cw[767] ^ cw[769] ^ cw[771] ^ cw[773] ^ cw[775] ^ cw[777] ^ cw[778] ^ cw[781] ^ cw[783] ^ cw[785] ^ cw[787] ^ cw[788] ^ cw[790] ^ cw[792] ^ cw[794] ^ cw[797] ^ cw[799] ^ cw[801] ^ cw[803] ^ cw[805] ^ cw[807] ^ cw[808] ^ cw[810] ^ cw[812] ^ cw[814] ^ cw[817] ^ cw[819] ^ cw[821] ^ cw[823] ^ cw[825] ^ cw[827] ^ cw[828] ^ cw[830] ^ cw[832] ^ cw[834] ^ cw[836] ^ cw[838] ^ cw[841] ^ cw[843] ^ cw[845] ^ cw[847] ^ cw[849] ^ cw[850] ^ cw[853] ^ cw[855] ^ cw[857] ^ cw[859] ^ cw[860] ^ cw[863] ^ cw[865] ^ cw[867] ^ cw[869] ^ cw[870] ^ cw[872] ^ cw[874] ^ cw[876] ^ cw[879] ^ cw[881] ^ cw[883] ^ cw[885] ^ cw[887] ^ cw[889] ^ cw[890] ^ cw[893] ^ cw[895] ^ cw[897] ^ cw[899] ^ cw[900] ^ cw[902] ^ cw[904] ^ cw[906] ^ cw[909] ^ cw[911] ^ cw[913] ^ cw[915] ^ cw[917] ^ cw[919] ^ cw[920] ^ cw[922] ^ cw[924] ^ cw[926] ^ cw[929] ^ cw[931] ^ cw[933] ^ cw[935] ^ cw[937] ^ cw[939] ^ cw[940] ^ cw[942] ^ cw[944] ^ cw[946] ^ cw[948] ^ cw[950] ^ cw[953] ^ cw[955] ^ cw[957] ^ cw[959] ^ cw[960] ^ cw[963] ^ cw[965] ^ cw[967] ^ cw[969] ^ cw[970] ^ cw[972] ^ cw[974] ^ cw[976] ^ cw[979] ^ cw[981] ^ cw[983] ^ cw[985] ^ cw[987] ^ cw[989] ^ cw[990] ^ cw[992] ^ cw[994] ^ cw[996] ^ cw[999] ^ cw[1001] ^ cw[1003] ^ cw[1005] ^ cw[1007] ^ cw[1009] ^ cw[1010] ^ cw[1012] ^ cw[1014] ^ cw[1016] ^ cw[1018] ^ cw[1020] ^ cw[1023] ^ cw[1025] ^ cw[1027] ^ cw[1029] ^ cw[1030] ^ cw[1032] ^ cw[1034] ^ cw[1036] ^ cw[1039] ^ cw[1041] ^ cw[1043] ^ cw[1045] ^ cw[1047] ^ cw[1049] ^ cw[1050] ^ cw[1052] ^ cw[1054] ^ cw[1056] ^ cw[1058] ^ cw[1060] ^ cw[1063] ^ cw[1065] ^ cw[1067] ^ cw[1069] ^ cw[1070] ^ cw[1072] ^ cw[1074] ^ cw[1076] ^ cw[1078] ^ cw[1080] ^ cw[1083] ^ cw[1085] ^ cw[1087] ^ cw[1089] ^ cw[1090] ^ cw[1092] ^ cw[1094] ^ cw[1096] ^ cw[1099] ^ cw[1101] ^ cw[1103] ^ cw[1104] ^ cw[1107] ^ cw[1109] ^ cw[1111] ^ cw[1113] ^ cw[1115] ^ cw[1116] ^ cw[1119] ^ cw[1121] ^ cw[1123] ^ cw[1125] ^ cw[1126] ^ cw[1129] ^ cw[1131] ^ cw[1133] ^ cw[1135] ^ cw[1136] ^ cw[1138] ^ cw[1140] ^ cw[1142] ^ cw[1145] ^ cw[1147] ^ cw[1149] ^ cw[1151] ^ cw[1153] ^ cw[1155] ^ cw[1157] ^ cw[1158] ^ cw[1161] ^ cw[1163] ^ cw[1165] ^ cw[1167] ^ cw[1168] ^ cw[1171] ^ cw[1173] ^ cw[1175] ^ cw[1177] ^ cw[1178] ^ cw[1180] ^ cw[1182] ^ cw[1184] ^ cw[1187] ^ cw[1189] ^ cw[1191] ^ cw[1193] ^ cw[1195] ^ cw[1197] ^ cw[1198] ^ cw[1201] ^ cw[1203] ^ cw[1205] ^ cw[1207] ^ cw[1208] ^ cw[1210] ^ cw[1212] ^ cw[1214] ^ cw[1217] ^ cw[1219] ^ cw[1221] ^ cw[1223] ^ cw[1225] ^ cw[1227] ^ cw[1228] ^ cw[1230] ^ cw[1232] ^ cw[1234] ^ cw[1237] ^ cw[1239] ^ cw[1241] ^ cw[1243] ^ cw[1245] ^ cw[1247] ^ cw[1248] ^ cw[1250] ^ cw[1252] ^ cw[1254] ^ cw[1256] ^ cw[1258] ^ cw[1261] ^ cw[1263] ^ cw[1265] ^ cw[1267] ^ cw[1269] ^ cw[1270] ^ cw[1273] ^ cw[1275] ^ cw[1277] ^ cw[1279] ^ cw[1280] ^ cw[1283] ^ cw[1285] ^ cw[1287] ^ cw[1289] ^ cw[1290] ^ cw[1292] ^ cw[1294] ^ cw[1296] ^ cw[1299] ^ cw[1301] ^ cw[1303] ^ cw[1305] ^ cw[1307] ^ cw[1309] ^ cw[1310] ^ cw[1313] ^ cw[1315] ^ cw[1317] ^ cw[1319] ^ cw[1320] ^ cw[1322] ^ cw[1324] ^ cw[1326] ^ cw[1329] ^ cw[1331] ^ cw[1333] ^ cw[1335] ^ cw[1337] ^ cw[1339] ^ cw[1340] ^ cw[1342] ^ cw[1344] ^ cw[1346] ^ cw[1349] ^ cw[1351] ^ cw[1353] ^ cw[1355] ^ cw[1357] ^ cw[1359] ^ cw[1360] ^ cw[1362] ^ cw[1364] ^ cw[1366] ^ cw[1368] ^ cw[1370] ^ cw[1373] ^ cw[1375] ^ cw[1377] ^ cw[1379] ^ cw[1380] ^ cw[1383] ^ cw[1385] ^ cw[1387] ^ cw[1389] ^ cw[1390] ^ cw[1392] ^ cw[1394] ^ cw[1396] ^ cw[1399] ^ cw[1401] ^ cw[1403] ^ cw[1405] ^ cw[1407] ^ cw[1409] ^ cw[1410] ^ cw[1412] ^ cw[1414] ^ cw[1416] ^ cw[1419] ^ cw[1421] ^ cw[1423] ^ cw[1425] ^ cw[1427] ^ cw[1429] ^ cw[1430] ^ cw[1432] ^ cw[1434] ^ cw[1436] ^ cw[1438] ^ cw[1440] ^ cw[1443] ^ cw[1445] ^ cw[1447] ^ cw[1449] ^ cw[1450] ^ cw[1452] ^ cw[1454] ^ cw[1456] ^ cw[1459] ^ cw[1461] ^ cw[1463] ^ cw[1465] ^ cw[1467] ^ cw[1469] ^ cw[1470] ^ cw[1472] ^ cw[1474] ^ cw[1476] ^ cw[1478] ^ cw[1480] ^ cw[1483] ^ cw[1485] ^ cw[1487] ^ cw[1489] ^ cw[1490] ^ cw[1492] ^ cw[1494] ^ cw[1496] ^ cw[1498] ^ cw[1500] ^ cw[1503] ^ cw[1505] ^ cw[1507] ^ cw[1509] ^ cw[1510] ^ cw[1512] ^ cw[1514] ^ cw[1516] ^ cw[1519] ^ cw[1521] ^ cw[1522] ^ cw[1525] ^ cw[1527] ^ cw[1529] ^ cw[1531] ^ cw[1532] ^ cw[1535] ^ cw[1537] ^ cw[1539] ^ cw[1541] ^ cw[1542] ^ cw[1544] ^ cw[1546] ^ cw[1548] ^ cw[1551] ^ cw[1553] ^ cw[1555] ^ cw[1557] ^ cw[1559] ^ cw[1561] ^ cw[1562] ^ cw[1565] ^ cw[1567] ^ cw[1569] ^ cw[1571] ^ cw[1572] ^ cw[1574] ^ cw[1576] ^ cw[1578] ^ cw[1581] ^ cw[1583] ^ cw[1585] ^ cw[1587] ^ cw[1589] ^ cw[1591] ^ cw[1592] ^ cw[1594] ^ cw[1596] ^ cw[1598] ^ cw[1601] ^ cw[1603] ^ cw[1605] ^ cw[1607] ^ cw[1609] ^ cw[1611] ^ cw[1612] ^ cw[1614] ^ cw[1616] ^ cw[1618] ^ cw[1620] ^ cw[1622] ^ cw[1625] ^ cw[1627] ^ cw[1629] ^ cw[1631] ^ cw[1632] ^ cw[1635] ^ cw[1637] ^ cw[1639] ^ cw[1641] ^ cw[1642] ^ cw[1644] ^ cw[1646] ^ cw[1648] ^ cw[1651] ^ cw[1653] ^ cw[1655] ^ cw[1657] ^ cw[1659] ^ cw[1661] ^ cw[1662] ^ cw[1664] ^ cw[1666] ^ cw[1668] ^ cw[1671] ^ cw[1673] ^ cw[1675] ^ cw[1677] ^ cw[1679] ^ cw[1681] ^ cw[1682] ^ cw[1684] ^ cw[1686] ^ cw[1688] ^ cw[1690] ^ cw[1692] ^ cw[1695] ^ cw[1697] ^ cw[1699] ^ cw[1701] ^ cw[1702] ^ cw[1704] ^ cw[1706] ^ cw[1708] ^ cw[1711] ^ cw[1713] ^ cw[1715] ^ cw[1717] ^ cw[1719] ^ cw[1721] ^ cw[1722] ^ cw[1724] ^ cw[1726] ^ cw[1728] ^ cw[1730] ^ cw[1732] ^ cw[1735] ^ cw[1737] ^ cw[1739] ^ cw[1741] ^ cw[1742] ^ cw[1744] ^ cw[1746] ^ cw[1748] ^ cw[1750] ^ cw[1752] ^ cw[1755] ^ cw[1757] ^ cw[1759] ^ cw[1761] ^ cw[1762] ^ cw[1764] ^ cw[1766] ^ cw[1768] ^ cw[1771] ^ cw[1772] ^ cw[1775] ^ cw[1777] ^ cw[1779] ^ cw[1781] ^ cw[1782] ^ cw[1784] ^ cw[1786] ^ cw[1788] ^ cw[1791] ^ cw[1793] ^ cw[1795] ^ cw[1797] ^ cw[1799] ^ cw[1801] ^ cw[1802] ^ cw[1804] ^ cw[1806] ^ cw[1808] ^ cw[1811] ^ cw[1813] ^ cw[1815] ^ cw[1817] ^ cw[1819] ^ cw[1821] ^ cw[1822] ^ cw[1824] ^ cw[1826] ^ cw[1828] ^ cw[1830] ^ cw[1832] ^ cw[1835] ^ cw[1837] ^ cw[1839] ^ cw[1841] ^ cw[1842] ^ cw[1844] ^ cw[1846] ^ cw[1848] ^ cw[1851] ^ cw[1853] ^ cw[1855] ^ cw[1857] ^ cw[1859] ^ cw[1861] ^ cw[1862] ^ cw[1864] ^ cw[1866] ^ cw[1868] ^ cw[1870] ^ cw[1872] ^ cw[1875] ^ cw[1877] ^ cw[1879] ^ cw[1881] ^ cw[1882] ^ cw[1884] ^ cw[1886] ^ cw[1888] ^ cw[1890] ^ cw[1892] ^ cw[1895] ^ cw[1897] ^ cw[1899] ^ cw[1901] ^ cw[1902] ^ cw[1904] ^ cw[1906] ^ cw[1908] ^ cw[1911] ^ cw[1912] ^ cw[1914] ^ cw[1916] ^ cw[1918] ^ cw[1921] ^ cw[1923] ^ cw[1925] ^ cw[1927] ^ cw[1929] ^ cw[1931] ^ cw[1932] ^ cw[1934] ^ cw[1936] ^ cw[1938] ^ cw[1940] ^ cw[1942] ^ cw[1945] ^ cw[1947] ^ cw[1949] ^ cw[1951] ^ cw[1952] ^ cw[1954] ^ cw[1956] ^ cw[1958] ^ cw[1960] ^ cw[1962] ^ cw[1965] ^ cw[1967] ^ cw[1969] ^ cw[1971] ^ cw[1972] ^ cw[1974] ^ cw[1976] ^ cw[1978] ^ cw[1981] ^ cw[1982] ^ cw[1984] ^ cw[1986] ^ cw[1988] ^ cw[1990] ^ cw[1992] ^ cw[1995] ^ cw[1997] ^ cw[1999] ^ cw[2001] ^ cw[2002] ^ cw[2004] ^ cw[2006] ^ cw[2008] ^ cw[2011] ^ cw[2012] ^ cw[2014] ^ cw[2016] ^ cw[2018] ^ cw[2021] ^ cw[2022] ^ cw[2024] ^ cw[2025] ^ cw[2026] ^ cw[2027] ^ cw[2029] ^ cw[2030] ^ cw[2031] ^ cw[2032] ^ cw[2033] ^ cw[2034] ^ cw[2035] ^ cw[2040];
    assign syndrome[6] = cw[1] ^ cw[3] ^ cw[5] ^ cw[7] ^ cw[8] ^ cw[11] ^ cw[13] ^ cw[15] ^ cw[17] ^ cw[19] ^ cw[21] ^ cw[23] ^ cw[25] ^ cw[26] ^ cw[29] ^ cw[31] ^ cw[33] ^ cw[35] ^ cw[37] ^ cw[39] ^ cw[41] ^ cw[42] ^ cw[45] ^ cw[47] ^ cw[49] ^ cw[51] ^ cw[53] ^ cw[55] ^ cw[56] ^ cw[59] ^ cw[61] ^ cw[63] ^ cw[65] ^ cw[67] ^ cw[68] ^ cw[71] ^ cw[73] ^ cw[75] ^ cw[77] ^ cw[79] ^ cw[80] ^ cw[82] ^ cw[84] ^ cw[86] ^ cw[88] ^ cw[91] ^ cw[93] ^ cw[95] ^ cw[97] ^ cw[99] ^ cw[101] ^ cw[103] ^ cw[105] ^ cw[107] ^ cw[109] ^ cw[111] ^ cw[113] ^ cw[115] ^ cw[116] ^ cw[119] ^ cw[121] ^ cw[123] ^ cw[125] ^ cw[127] ^ cw[129] ^ cw[131] ^ cw[132] ^ cw[135] ^ cw[137] ^ cw[139] ^ cw[141] ^ cw[143] ^ cw[145] ^ cw[146] ^ cw[149] ^ cw[151] ^ cw[153] ^ cw[155] ^ cw[157] ^ cw[158] ^ cw[161] ^ cw[163] ^ cw[165] ^ cw[167] ^ cw[169] ^ cw[170] ^ cw[172] ^ cw[174] ^ cw[176] ^ cw[178] ^ cw[181] ^ cw[183] ^ cw[185] ^ cw[187] ^ cw[189] ^ cw[191] ^ cw[193] ^ cw[195] ^ cw[197] ^ cw[199] ^ cw[201] ^ cw[203] ^ cw[204] ^ cw[207] ^ cw[209] ^ cw[211] ^ cw[213] ^ cw[215] ^ cw[217] ^ cw[218] ^ cw[221] ^ cw[223] ^ cw[225] ^ cw[227] ^ cw[229] ^ cw[230] ^ cw[233] ^ cw[235] ^ cw[237] ^ cw[239] ^ cw[241] ^ cw[242] ^ cw[244] ^ cw[246] ^ cw[248] ^ cw[250] ^ cw[253] ^ cw[255] ^ cw[257] ^ cw[259] ^ cw[261] ^ cw[263] ^ cw[265] ^ cw[267] ^ cw[269] ^ cw[271] ^ cw[273] ^ cw[274] ^ cw[277] ^ cw[279] ^ cw[281] ^ cw[283] ^ cw[285] ^ cw[286] ^ cw[289] ^ cw[291] ^ cw[293] ^ cw[295] ^ cw[297] ^ cw[298] ^ cw[300] ^ cw[302] ^ cw[304] ^ cw[306] ^ cw[309] ^ cw[311] ^ cw[313] ^ cw[315] ^ cw[317] ^ cw[319] ^ cw[321] ^ cw[323] ^ cw[325] ^ cw[327] ^ cw[328] ^ cw[331] ^ cw[333] ^ cw[335] ^ cw[337] ^ cw[339] ^ cw[340] ^ cw[342] ^ cw[344] ^ cw[346] ^ cw[348] ^ cw[351] ^ cw[353] ^ cw[355] ^ cw[357] ^ cw[359] ^ cw[361] ^ cw[363] ^ cw[365] ^ cw[367] ^ cw[369] ^ cw[370] ^ cw[372] ^ cw[374] ^ cw[376] ^ cw[378] ^ cw[381] ^ cw[383] ^ cw[385] ^ cw[387] ^ cw[389] ^ cw[391] ^ cw[393] ^ cw[395] ^ cw[397] ^ cw[399] ^ cw[400] ^ cw[402] ^ cw[404] ^ cw[406] ^ cw[408] ^ cw[410] ^ cw[412] ^ cw[414] ^ cw[416] ^ cw[418] ^ cw[421] ^ cw[423] ^ cw[425] ^ cw[427] ^ cw[429] ^ cw[431] ^ cw[433] ^ cw[435] ^ cw[437] ^ cw[439] ^ cw[441] ^ cw[443] ^ cw[444] ^ cw[447] ^ cw[449] ^ cw[451] ^ cw[453] ^ cw[455] ^ cw[457] ^ cw[458] ^ cw[461] ^ cw[463] ^ cw[465] ^ cw[467] ^ cw[469] ^ cw[470] ^ cw[473] ^ cw[475] ^ cw[477] ^ cw[479] ^ cw[481] ^ cw[482] ^ cw[484] ^ cw[486] ^ cw[488] ^ cw[490] ^ cw[493] ^ cw[495] ^ cw[497] ^ cw[499] ^ cw[501] ^ cw[503] ^ cw[505] ^ cw[507] ^ cw[509] ^ cw[511] ^ cw[513] ^ cw[514] ^ cw[517] ^ cw[519] ^ cw[521] ^ cw[523] ^ cw[525] ^ cw[526] ^ cw[529] ^ cw[531] ^ cw[533] ^ cw[535] ^ cw[537] ^ cw[538] ^ cw[540] ^ cw[542] ^ cw[544] ^ cw[546] ^ cw[549] ^ cw[551] ^ cw[553] ^ cw[555] ^ cw[557] ^ cw[559] ^ cw[561] ^ cw[563] ^ cw[565] ^ cw[567] ^ cw[568] ^ cw[571] ^ cw[573] ^ cw[575] ^ cw[577] ^ cw[579] ^ cw[580] ^ cw[582] ^ cw[584] ^ cw[586] ^ cw[588] ^ cw[591] ^ cw[593] ^ cw[595] ^ cw[597] ^ cw[599] ^ cw[601] ^ cw[603] ^ cw[605] ^ cw[607] ^ cw[609] ^ cw[610] ^ cw[612] ^ cw[614] ^ cw[616] ^ cw[618] ^ cw[621] ^ cw[623] ^ cw[625] ^ cw[627] ^ cw[629] ^ cw[631] ^ cw[633] ^ cw[635] ^ cw[637] ^ cw[639] ^ cw[640] ^ cw[642] ^ cw[644] ^ cw[646] ^ cw[648] ^ cw[650] ^ cw[652] ^ cw[654] ^ cw[656] ^ cw[658] ^ cw[661] ^ cw[663] ^ cw[665] ^ cw[667] ^ cw[669] ^ cw[671] ^ cw[673] ^ cw[675] ^ cw[677] ^ cw[679] ^ cw[681] ^ cw[682] ^ cw[685] ^ cw[687] ^ cw[689] ^ cw[691] ^ cw[693] ^ cw[694] ^ cw[697] ^ cw[699] ^ cw[701] ^ cw[703] ^ cw[705] ^ cw[706] ^ cw[708] ^ cw[710] ^ cw[712] ^ cw[714] ^ cw[717] ^ cw[719] ^ cw[721] ^ cw[723] ^ cw[725] ^ cw[727] ^ cw[729] ^ cw[731] ^ cw[733] ^ cw[735] ^ cw[736] ^ cw[739] ^ cw[741] ^ cw[743] ^ cw[745] ^ cw[747] ^ cw[748] ^ cw[750] ^ cw[752] ^ cw[754] ^ cw[756] ^ cw[759] ^ cw[761] ^ cw[763] ^ cw[765] ^ cw[767] ^ cw[769] ^ cw[771] ^ cw[773] ^ cw[775] ^ cw[777] ^ cw[778] ^ cw[780] ^ cw[782] ^ cw[784] ^ cw[786] ^ cw[789] ^ cw[791] ^ cw[793] ^ cw[795] ^ cw[797] ^ cw[799] ^ cw[801] ^ cw[803] ^ cw[805] ^ cw[807] ^ cw[808] ^ cw[810] ^ cw[812] ^ cw[814] ^ cw[816] ^ cw[818] ^ cw[820] ^ cw[822] ^ cw[824] ^ cw[826] ^ cw[829] ^ cw[831] ^ cw[833] ^ cw[835] ^ cw[837] ^ cw[839] ^ cw[841] ^ cw[843] ^ cw[845] ^ cw[847] ^ cw[848] ^ cw[851] ^ cw[853] ^ cw[855] ^ cw[857] ^ cw[859] ^ cw[860] ^ cw[862] ^ cw[864] ^ cw[866] ^ cw[868] ^ cw[871] ^ cw[873] ^ cw[875] ^ cw[877] ^ cw[879] ^ cw[881] ^ cw[883] ^ cw[885] ^ cw[887] ^ cw[889] ^ cw[890] ^ cw[892] ^ cw[894] ^ cw[896] ^ cw[898] ^ cw[901] ^ cw[903] ^ cw[905] ^ cw[907] ^ cw[909] ^ cw[911] ^ cw[913] ^ cw[915] ^ cw[917] ^ cw[919] ^ cw[920] ^ cw[922] ^ cw[924] ^ cw[926] ^ cw[928] ^ cw[930] ^ cw[932] ^ cw[934] ^ cw[936] ^ cw[938] ^ cw[941] ^ cw[943] ^ cw[945] ^ cw[947] ^ cw[949] ^ cw[951] ^ cw[953] ^ cw[955] ^ cw[957] ^ cw[959] ^ cw[960] ^ cw[962] ^ cw[964] ^ cw[966] ^ cw[968] ^ cw[971] ^ cw[973] ^ cw[975] ^ cw[977] ^ cw[979] ^ cw[981] ^ cw[983] ^ cw[985] ^ cw[987] ^ cw[989] ^ cw[990] ^ cw[992] ^ cw[994] ^ cw[996] ^ cw[998] ^ cw[1000] ^ cw[1002] ^ cw[1004] ^ cw[1006] ^ cw[1008] ^ cw[1011] ^ cw[1013] ^ cw[1015] ^ cw[1017] ^ cw[1019] ^ cw[1021] ^ cw[1023] ^ cw[1025] ^ cw[1027] ^ cw[1029] ^ cw[1030] ^ cw[1032] ^ cw[1034] ^ cw[1036] ^ cw[1038] ^ cw[1040] ^ cw[1042] ^ cw[1044] ^ cw[1046] ^ cw[1048] ^ cw[1051] ^ cw[1053] ^ cw[1055] ^ cw[1057] ^ cw[1059] ^ cw[1061] ^ cw[1063] ^ cw[1065] ^ cw[1067] ^ cw[1069] ^ cw[1070] ^ cw[1072] ^ cw[1074] ^ cw[1076] ^ cw[1078] ^ cw[1080] ^ cw[1082] ^ cw[1084] ^ cw[1086] ^ cw[1088] ^ cw[1091] ^ cw[1093] ^ cw[1095] ^ cw[1097] ^ cw[1099] ^ cw[1101] ^ cw[1102] ^ cw[1105] ^ cw[1107] ^ cw[1109] ^ cw[1111] ^ cw[1113] ^ cw[1114] ^ cw[1117] ^ cw[1119] ^ cw[1121] ^ cw[1123] ^ cw[1125] ^ cw[1126] ^ cw[1128] ^ cw[1130] ^ cw[1132] ^ cw[1134] ^ cw[1137] ^ cw[1139] ^ cw[1141] ^ cw[1143] ^ cw[1145] ^ cw[1147] ^ cw[1149] ^ cw[1151] ^ cw[1153] ^ cw[1155] ^ cw[1156] ^ cw[1159] ^ cw[1161] ^ cw[1163] ^ cw[1165] ^ cw[1167] ^ cw[1168] ^ cw[1170] ^ cw[1172] ^ cw[1174] ^ cw[1176] ^ cw[1179] ^ cw[1181] ^ cw[1183] ^ cw[1185] ^ cw[1187] ^ cw[1189] ^ cw[1191] ^ cw[1193] ^ cw[1195] ^ cw[1197] ^ cw[1198] ^ cw[1200] ^ cw[1202] ^ cw[1204] ^ cw[1206] ^ cw[1209] ^ cw[1211] ^ cw[1213] ^ cw[1215] ^ cw[1217] ^ cw[1219] ^ cw[1221] ^ cw[1223] ^ cw[1225] ^ cw[1227] ^ cw[1228] ^ cw[1230] ^ cw[1232] ^ cw[1234] ^ cw[1236] ^ cw[1238] ^ cw[1240] ^ cw[1242] ^ cw[1244] ^ cw[1246] ^ cw[1249] ^ cw[1251] ^ cw[1253] ^ cw[1255] ^ cw[1257] ^ cw[1259] ^ cw[1261] ^ cw[1263] ^ cw[1265] ^ cw[1267] ^ cw[1268] ^ cw[1271] ^ cw[1273] ^ cw[1275] ^ cw[1277] ^ cw[1279] ^ cw[1280] ^ cw[1282] ^ cw[1284] ^ cw[1286] ^ cw[1288] ^ cw[1291] ^ cw[1293] ^ cw[1295] ^ cw[1297] ^ cw[1299] ^ cw[1301] ^ cw[1303] ^ cw[1305] ^ cw[1307] ^ cw[1309] ^ cw[1310] ^ cw[1312] ^ cw[1314] ^ cw[1316] ^ cw[1318] ^ cw[1321] ^ cw[1323] ^ cw[1325] ^ cw[1327] ^ cw[1329] ^ cw[1331] ^ cw[1333] ^ cw[1335] ^ cw[1337] ^ cw[1339] ^ cw[1340] ^ cw[1342] ^ cw[1344] ^ cw[1346] ^ cw[1348] ^ cw[1350] ^ cw[1352] ^ cw[1354] ^ cw[1356] ^ cw[1358] ^ cw[1361] ^ cw[1363] ^ cw[1365] ^ cw[1367] ^ cw[1369] ^ cw[1371] ^ cw[1373] ^ cw[1375] ^ cw[1377] ^ cw[1379] ^ cw[1380] ^ cw[1382] ^ cw[1384] ^ cw[1386] ^ cw[1388] ^ cw[1391] ^ cw[1393] ^ cw[1395] ^ cw[1397] ^ cw[1399] ^ cw[1401] ^ cw[1403] ^ cw[1405] ^ cw[1407] ^ cw[1409] ^ cw[1410] ^ cw[1412] ^ cw[1414] ^ cw[1416] ^ cw[1418] ^ cw[1420] ^ cw[1422] ^ cw[1424] ^ cw[1426] ^ cw[1428] ^ cw[1431] ^ cw[1433] ^ cw[1435] ^ cw[1437] ^ cw[1439] ^ cw[1441] ^ cw[1443] ^ cw[1445] ^ cw[1447] ^ cw[1449] ^ cw[1450] ^ cw[1452] ^ cw[1454] ^ cw[1456] ^ cw[1458] ^ cw[1460] ^ cw[1462] ^ cw[1464] ^ cw[1466] ^ cw[1468] ^ cw[1471] ^ cw[1473] ^ cw[1475] ^ cw[1477] ^ cw[1479] ^ cw[1481] ^ cw[1483] ^ cw[1485] ^ cw[1487] ^ cw[1489] ^ cw[1490] ^ cw[1492] ^ cw[1494] ^ cw[1496] ^ cw[1498] ^ cw[1500] ^ cw[1502] ^ cw[1504] ^ cw[1506] ^ cw[1508] ^ cw[1511] ^ cw[1513] ^ cw[1515] ^ cw[1517] ^ cw[1519] ^ cw[1520] ^ cw[1523] ^ cw[1525] ^ cw[1527] ^ cw[1529] ^ cw[1531] ^ cw[1532] ^ cw[1534] ^ cw[1536] ^ cw[1538] ^ cw[1540] ^ cw[1543] ^ cw[1545] ^ cw[1547] ^ cw[1549] ^ cw[1551] ^ cw[1553] ^ cw[1555] ^ cw[1557] ^ cw[1559] ^ cw[1561] ^ cw[1562] ^ cw[1564] ^ cw[1566] ^ cw[1568] ^ cw[1570] ^ cw[1573] ^ cw[1575] ^ cw[1577] ^ cw[1579] ^ cw[1581] ^ cw[1583] ^ cw[1585] ^ cw[1587] ^ cw[1589] ^ cw[1591] ^ cw[1592] ^ cw[1594] ^ cw[1596] ^ cw[1598] ^ cw[1600] ^ cw[1602] ^ cw[1604] ^ cw[1606] ^ cw[1608] ^ cw[1610] ^ cw[1613] ^ cw[1615] ^ cw[1617] ^ cw[1619] ^ cw[1621] ^ cw[1623] ^ cw[1625] ^ cw[1627] ^ cw[1629] ^ cw[1631] ^ cw[1632] ^ cw[1634] ^ cw[1636] ^ cw[1638] ^ cw[1640] ^ cw[1643] ^ cw[1645] ^ cw[1647] ^ cw[1649] ^ cw[1651] ^ cw[1653] ^ cw[1655] ^ cw[1657] ^ cw[1659] ^ cw[1661] ^ cw[1662] ^ cw[1664] ^ cw[1666] ^ cw[1668] ^ cw[1670] ^ cw[1672] ^ cw[1674] ^ cw[1676] ^ cw[1678] ^ cw[1680] ^ cw[1683] ^ cw[1685] ^ cw[1687] ^ cw[1689] ^ cw[1691] ^ cw[1693] ^ cw[1695] ^ cw[1697] ^ cw[1699] ^ cw[1701] ^ cw[1702] ^ cw[1704] ^ cw[1706] ^ cw[1708] ^ cw[1710] ^ cw[1712] ^ cw[1714] ^ cw[1716] ^ cw[1718] ^ cw[1720] ^ cw[1723] ^ cw[1725] ^ cw[1727] ^ cw[1729] ^ cw[1731] ^ cw[1733] ^ cw[1735] ^ cw[1737] ^ cw[1739] ^ cw[1741] ^ cw[1742] ^ cw[1744] ^ cw[1746] ^ cw[1748] ^ cw[1750] ^ cw[1752] ^ cw[1754] ^ cw[1756] ^ cw[1758] ^ cw[1760] ^ cw[1763] ^ cw[1765] ^ cw[1767] ^ cw[1769] ^ cw[1771] ^ cw[1772] ^ cw[1774] ^ cw[1776] ^ cw[1778] ^ cw[1780] ^ cw[1783] ^ cw[1785] ^ cw[1787] ^ cw[1789] ^ cw[1791] ^ cw[1793] ^ cw[1795] ^ cw[1797] ^ cw[1799] ^ cw[1801] ^ cw[1802] ^ cw[1804] ^ cw[1806] ^ cw[1808] ^ cw[1810] ^ cw[1812] ^ cw[1814] ^ cw[1816] ^ cw[1818] ^ cw[1820] ^ cw[1823] ^ cw[1825] ^ cw[1827] ^ cw[1829] ^ cw[1831] ^ cw[1833] ^ cw[1835] ^ cw[1837] ^ cw[1839] ^ cw[1841] ^ cw[1842] ^ cw[1844] ^ cw[1846] ^ cw[1848] ^ cw[1850] ^ cw[1852] ^ cw[1854] ^ cw[1856] ^ cw[1858] ^ cw[1860] ^ cw[1863] ^ cw[1865] ^ cw[1867] ^ cw[1869] ^ cw[1871] ^ cw[1873] ^ cw[1875] ^ cw[1877] ^ cw[1879] ^ cw[1881] ^ cw[1882] ^ cw[1884] ^ cw[1886] ^ cw[1888] ^ cw[1890] ^ cw[1892] ^ cw[1894] ^ cw[1896] ^ cw[1898] ^ cw[1900] ^ cw[1903] ^ cw[1905] ^ cw[1907] ^ cw[1909] ^ cw[1911] ^ cw[1912] ^ cw[1914] ^ cw[1916] ^ cw[1918] ^ cw[1920] ^ cw[1922] ^ cw[1924] ^ cw[1926] ^ cw[1928] ^ cw[1930] ^ cw[1933] ^ cw[1935] ^ cw[1937] ^ cw[1939] ^ cw[1941] ^ cw[1943] ^ cw[1945] ^ cw[1947] ^ cw[1949] ^ cw[1951] ^ cw[1952] ^ cw[1954] ^ cw[1956] ^ cw[1958] ^ cw[1960] ^ cw[1962] ^ cw[1964] ^ cw[1966] ^ cw[1968] ^ cw[1970] ^ cw[1973] ^ cw[1975] ^ cw[1977] ^ cw[1979] ^ cw[1981] ^ cw[1982] ^ cw[1984] ^ cw[1986] ^ cw[1988] ^ cw[1990] ^ cw[1992] ^ cw[1994] ^ cw[1996] ^ cw[1998] ^ cw[2000] ^ cw[2003] ^ cw[2005] ^ cw[2007] ^ cw[2009] ^ cw[2011] ^ cw[2012] ^ cw[2014] ^ cw[2016] ^ cw[2018] ^ cw[2020] ^ cw[2023] ^ cw[2024] ^ cw[2025] ^ cw[2026] ^ cw[2027] ^ cw[2028] ^ cw[2030] ^ cw[2031] ^ cw[2032] ^ cw[2033] ^ cw[2034] ^ cw[2035] ^ cw[2041];
    assign syndrome[5] = cw[1] ^ cw[3] ^ cw[5] ^ cw[6] ^ cw[9] ^ cw[11] ^ cw[13] ^ cw[15] ^ cw[17] ^ cw[19] ^ cw[21] ^ cw[23] ^ cw[24] ^ cw[27] ^ cw[29] ^ cw[31] ^ cw[33] ^ cw[35] ^ cw[37] ^ cw[39] ^ cw[40] ^ cw[43] ^ cw[45] ^ cw[47] ^ cw[49] ^ cw[51] ^ cw[53] ^ cw[54] ^ cw[57] ^ cw[59] ^ cw[61] ^ cw[63] ^ cw[65] ^ cw[67] ^ cw[68] ^ cw[70] ^ cw[72] ^ cw[74] ^ cw[76] ^ cw[78] ^ cw[81] ^ cw[83] ^ cw[85] ^ cw[87] ^ cw[89] ^ cw[91] ^ cw[93] ^ cw[95] ^ cw[97] ^ cw[99] ^ cw[101] ^ cw[103] ^ cw[105] ^ cw[107] ^ cw[109] ^ cw[111] ^ cw[113] ^ cw[114] ^ cw[117] ^ cw[119] ^ cw[121] ^ cw[123] ^ cw[125] ^ cw[127] ^ cw[129] ^ cw[130] ^ cw[133] ^ cw[135] ^ cw[137] ^ cw[139] ^ cw[141] ^ cw[143] ^ cw[144] ^ cw[147] ^ cw[149] ^ cw[151] ^ cw[153] ^ cw[155] ^ cw[157] ^ cw[158] ^ cw[160] ^ cw[162] ^ cw[164] ^ cw[166] ^ cw[168] ^ cw[171] ^ cw[173] ^ cw[175] ^ cw[177] ^ cw[179] ^ cw[181] ^ cw[183] ^ cw[185] ^ cw[187] ^ cw[189] ^ cw[191] ^ cw[193] ^ cw[195] ^ cw[197] ^ cw[199] ^ cw[201] ^ cw[202] ^ cw[205] ^ cw[207] ^ cw[209] ^ cw[211] ^ cw[213] ^ cw[215] ^ cw[216] ^ cw[219] ^ cw[221] ^ cw[223] ^ cw[225] ^ cw[227] ^ cw[229] ^ cw[230] ^ cw[232] ^ cw[234] ^ cw[236] ^ cw[238] ^ cw[240] ^ cw[243] ^ cw[245] ^ cw[247] ^ cw[249] ^ cw[251] ^ cw[253] ^ cw[255] ^ cw[257] ^ cw[259] ^ cw[261] ^ cw[263] ^ cw[265] ^ cw[267] ^ cw[269] ^ cw[271] ^ cw[272] ^ cw[275] ^ cw[277] ^ cw[279] ^ cw[281] ^ cw[283] ^ cw[285] ^ cw[286] ^ cw[288] ^ cw[290] ^ cw[292] ^ cw[294] ^ cw[296] ^ cw[299] ^ cw[301] ^ cw[303] ^ cw[305] ^ cw[307] ^ cw[309] ^ cw[311] ^ cw[313] ^ cw[315] ^ cw[317] ^ cw[319] ^ cw[321] ^ cw[323] ^ cw[325] ^ cw[327] ^ cw[328] ^ cw[330] ^ cw[332] ^ cw[334] ^ cw[336] ^ cw[338] ^ cw[341] ^ cw[343] ^ cw[345] ^ cw[347] ^ cw[349] ^ cw[351] ^ cw[353] ^ cw[355] ^ cw[357] ^ cw[359] ^ cw[361] ^ cw[363] ^ cw[365] ^ cw[367] ^ cw[369] ^ cw[370] ^ cw[372] ^ cw[374] ^ cw[376] ^ cw[378] ^ cw[380] ^ cw[382] ^ cw[384] ^ cw[386] ^ cw[388] ^ cw[390] ^ cw[392] ^ cw[394] ^ cw[396] ^ cw[398] ^ cw[401] ^ cw[403] ^ cw[405] ^ cw[407] ^ cw[409] ^ cw[411] ^ cw[413] ^ cw[415] ^ cw[417] ^ cw[419] ^ cw[421] ^ cw[423] ^ cw[425] ^ cw[427] ^ cw[429] ^ cw[431] ^ cw[433] ^ cw[435] ^ cw[437] ^ cw[439] ^ cw[441] ^ cw[442] ^ cw[445] ^ cw[447] ^ cw[449] ^ cw[451] ^ cw[453] ^ cw[455] ^ cw[456] ^ cw[459] ^ cw[461] ^ cw[463] ^ cw[465] ^ cw[467] ^ cw[469] ^ cw[470] ^ cw[472] ^ cw[474] ^ cw[476] ^ cw[478] ^ cw[480] ^ cw[483] ^ cw[485] ^ cw[487] ^ cw[489] ^ cw[491] ^ cw[493] ^ cw[495] ^ cw[497] ^ cw[499] ^ cw[501] ^ cw[503] ^ cw[505] ^ cw[507] ^ cw[509] ^ cw[511] ^ cw[512] ^ cw[515] ^ cw[517] ^ cw[519] ^ cw[521] ^ cw[523] ^ cw[525] ^ cw[526] ^ cw[528] ^ cw[530] ^ cw[532] ^ cw[534] ^ cw[536] ^ cw[539] ^ cw[541] ^ cw[543] ^ cw[545] ^ cw[547] ^ cw[549] ^ cw[551] ^ cw[553] ^ cw[555] ^ cw[557] ^ cw[559] ^ cw[561] ^ cw[563] ^ cw[565] ^ cw[567] ^ cw[568] ^ cw[570] ^ cw[572] ^ cw[574] ^ cw[576] ^ cw[578] ^ cw[581] ^ cw[583] ^ cw[585] ^ cw[587] ^ cw[589] ^ cw[591] ^ cw[593] ^ cw[595] ^ cw[597] ^ cw[599] ^ cw[601] ^ cw[603] ^ cw[605] ^ cw[607] ^ cw[609] ^ cw[610] ^ cw[612] ^ cw[614] ^ cw[616] ^ cw[618] ^ cw[620] ^ cw[622] ^ cw[624] ^ cw[626] ^ cw[628] ^ cw[630] ^ cw[632] ^ cw[634] ^ cw[636] ^ cw[638] ^ cw[641] ^ cw[643] ^ cw[645] ^ cw[647] ^ cw[649] ^ cw[651] ^ cw[653] ^ cw[655] ^ cw[657] ^ cw[659] ^ cw[661] ^ cw[663] ^ cw[665] ^ cw[667] ^ cw[669] ^ cw[671] ^ cw[673] ^ cw[675] ^ cw[677] ^ cw[679] ^ cw[680] ^ cw[683] ^ cw[685] ^ cw[687] ^ cw[689] ^ cw[691] ^ cw[693] ^ cw[694] ^ cw[696] ^ cw[698] ^ cw[700] ^ cw[702] ^ cw[704] ^ cw[707] ^ cw[709] ^ cw[711] ^ cw[713] ^ cw[715] ^ cw[717] ^ cw[719] ^ cw[721] ^ cw[723] ^ cw[725] ^ cw[727] ^ cw[729] ^ cw[731] ^ cw[733] ^ cw[735] ^ cw[736] ^ cw[738] ^ cw[740] ^ cw[742] ^ cw[744] ^ cw[746] ^ cw[749] ^ cw[751] ^ cw[753] ^ cw[755] ^ cw[757] ^ cw[759] ^ cw[761] ^ cw[763] ^ cw[765] ^ cw[767] ^ cw[769] ^ cw[771] ^ cw[773] ^ cw[775] ^ cw[777] ^ cw[778] ^ cw[780] ^ cw[782] ^ cw[784] ^ cw[786] ^ cw[788] ^ cw[790] ^ cw[792] ^ cw[794] ^ cw[796] ^ cw[798] ^ cw[800] ^ cw[802] ^ cw[804] ^ cw[806] ^ cw[809] ^ cw[811] ^ cw[813] ^ cw[815] ^ cw[817] ^ cw[819] ^ cw[821] ^ cw[823] ^ cw[825] ^ cw[827] ^ cw[829] ^ cw[831] ^ cw[833] ^ cw[835] ^ cw[837] ^ cw[839] ^ cw[841] ^ cw[843] ^ cw[845] ^ cw[847] ^ cw[848] ^ cw[850] ^ cw[852] ^ cw[854] ^ cw[856] ^ cw[858] ^ cw[861] ^ cw[863] ^ cw[865] ^ cw[867] ^ cw[869] ^ cw[871] ^ cw[873] ^ cw[875] ^ cw[877] ^ cw[879] ^ cw[881] ^ cw[883] ^ cw[885] ^ cw[887] ^ cw[889] ^ cw[890] ^ cw[892] ^ cw[894] ^ cw[896] ^ cw[898] ^ cw[900] ^ cw[902] ^ cw[904] ^ cw[906] ^ cw[908] ^ cw[910] ^ cw[912] ^ cw[914] ^ cw[916] ^ cw[918] ^ cw[921] ^ cw[923] ^ cw[925] ^ cw[927] ^ cw[929] ^ cw[931] ^ cw[933] ^ cw[935] ^ cw[937] ^ cw[939] ^ cw[941] ^ cw[943] ^ cw[945] ^ cw[947] ^ cw[949] ^ cw[951] ^ cw[953] ^ cw[955] ^ cw[957] ^ cw[959] ^ cw[960] ^ cw[962] ^ cw[964] ^ cw[966] ^ cw[968] ^ cw[970] ^ cw[972] ^ cw[974] ^ cw[976] ^ cw[978] ^ cw[980] ^ cw[982] ^ cw[984] ^ cw[986] ^ cw[988] ^ cw[991] ^ cw[993] ^ cw[995] ^ cw[997] ^ cw[999] ^ cw[1001] ^ cw[1003] ^ cw[1005] ^ cw[1007] ^ cw[1009] ^ cw[1011] ^ cw[1013] ^ cw[1015] ^ cw[1017] ^ cw[1019] ^ cw[1021] ^ cw[1023] ^ cw[1025] ^ cw[1027] ^ cw[1029] ^ cw[1030] ^ cw[1032] ^ cw[1034] ^ cw[1036] ^ cw[1038] ^ cw[1040] ^ cw[1042] ^ cw[1044] ^ cw[1046] ^ cw[1048] ^ cw[1050] ^ cw[1052] ^ cw[1054] ^ cw[1056] ^ cw[1058] ^ cw[1060] ^ cw[1062] ^ cw[1064] ^ cw[1066] ^ cw[1068] ^ cw[1071] ^ cw[1073] ^ cw[1075] ^ cw[1077] ^ cw[1079] ^ cw[1081] ^ cw[1083] ^ cw[1085] ^ cw[1087] ^ cw[1089] ^ cw[1091] ^ cw[1093] ^ cw[1095] ^ cw[1097] ^ cw[1099] ^ cw[1100] ^ cw[1103] ^ cw[1105] ^ cw[1107] ^ cw[1109] ^ cw[1111] ^ cw[1113] ^ cw[1114] ^ cw[1116] ^ cw[1118] ^ cw[1120] ^ cw[1122] ^ cw[1124] ^ cw[1127] ^ cw[1129] ^ cw[1131] ^ cw[1133] ^ cw[1135] ^ cw[1137] ^ cw[1139] ^ cw[1141] ^ cw[1143] ^ cw[1145] ^ cw[1147] ^ cw[1149] ^ cw[1151] ^ cw[1153] ^ cw[1155] ^ cw[1156] ^ cw[1158] ^ cw[1160] ^ cw[1162] ^ cw[1164] ^ cw[1166] ^ cw[1169] ^ cw[1171] ^ cw[1173] ^ cw[1175] ^ cw[1177] ^ cw[1179] ^ cw[1181] ^ cw[1183] ^ cw[1185] ^ cw[1187] ^ cw[1189] ^ cw[1191] ^ cw[1193] ^ cw[1195] ^ cw[1197] ^ cw[1198] ^ cw[1200] ^ cw[1202] ^ cw[1204] ^ cw[1206] ^ cw[1208] ^ cw[1210] ^ cw[1212] ^ cw[1214] ^ cw[1216] ^ cw[1218] ^ cw[1220] ^ cw[1222] ^ cw[1224] ^ cw[1226] ^ cw[1229] ^ cw[1231] ^ cw[1233] ^ cw[1235] ^ cw[1237] ^ cw[1239] ^ cw[1241] ^ cw[1243] ^ cw[1245] ^ cw[1247] ^ cw[1249] ^ cw[1251] ^ cw[1253] ^ cw[1255] ^ cw[1257] ^ cw[1259] ^ cw[1261] ^ cw[1263] ^ cw[1265] ^ cw[1267] ^ cw[1268] ^ cw[1270] ^ cw[1272] ^ cw[1274] ^ cw[1276] ^ cw[1278] ^ cw[1281] ^ cw[1283] ^ cw[1285] ^ cw[1287] ^ cw[1289] ^ cw[1291] ^ cw[1293] ^ cw[1295] ^ cw[1297] ^ cw[1299] ^ cw[1301] ^ cw[1303] ^ cw[1305] ^ cw[1307] ^ cw[1309] ^ cw[1310] ^ cw[1312] ^ cw[1314] ^ cw[1316] ^ cw[1318] ^ cw[1320] ^ cw[1322] ^ cw[1324] ^ cw[1326] ^ cw[1328] ^ cw[1330] ^ cw[1332] ^ cw[1334] ^ cw[1336] ^ cw[1338] ^ cw[1341] ^ cw[1343] ^ cw[1345] ^ cw[1347] ^ cw[1349] ^ cw[1351] ^ cw[1353] ^ cw[1355] ^ cw[1357] ^ cw[1359] ^ cw[1361] ^ cw[1363] ^ cw[1365] ^ cw[1367] ^ cw[1369] ^ cw[1371] ^ cw[1373] ^ cw[1375] ^ cw[1377] ^ cw[1379] ^ cw[1380] ^ cw[1382] ^ cw[1384] ^ cw[1386] ^ cw[1388] ^ cw[1390] ^ cw[1392] ^ cw[1394] ^ cw[1396] ^ cw[1398] ^ cw[1400] ^ cw[1402] ^ cw[1404] ^ cw[1406] ^ cw[1408] ^ cw[1411] ^ cw[1413] ^ cw[1415] ^ cw[1417] ^ cw[1419] ^ cw[1421] ^ cw[1423] ^ cw[1425] ^ cw[1427] ^ cw[1429] ^ cw[1431] ^ cw[1433] ^ cw[1435] ^ cw[1437] ^ cw[1439] ^ cw[1441] ^ cw[1443] ^ cw[1445] ^ cw[1447] ^ cw[1449] ^ cw[1450] ^ cw[1452] ^ cw[1454] ^ cw[1456] ^ cw[1458] ^ cw[1460] ^ cw[1462] ^ cw[1464] ^ cw[1466] ^ cw[1468] ^ cw[1470] ^ cw[1472] ^ cw[1474] ^ cw[1476] ^ cw[1478] ^ cw[1480] ^ cw[1482] ^ cw[1484] ^ cw[1486] ^ cw[1488] ^ cw[1491] ^ cw[1493] ^ cw[1495] ^ cw[1497] ^ cw[1499] ^ cw[1501] ^ cw[1503] ^ cw[1505] ^ cw[1507] ^ cw[1509] ^ cw[1511] ^ cw[1513] ^ cw[1515] ^ cw[1517] ^ cw[1519] ^ cw[1520] ^ cw[1522] ^ cw[1524] ^ cw[1526] ^ cw[1528] ^ cw[1530] ^ cw[1533] ^ cw[1535] ^ cw[1537] ^ cw[1539] ^ cw[1541] ^ cw[1543] ^ cw[1545] ^ cw[1547] ^ cw[1549] ^ cw[1551] ^ cw[1553] ^ cw[1555] ^ cw[1557] ^ cw[1559] ^ cw[1561] ^ cw[1562] ^ cw[1564] ^ cw[1566] ^ cw[1568] ^ cw[1570] ^ cw[1572] ^ cw[1574] ^ cw[1576] ^ cw[1578] ^ cw[1580] ^ cw[1582] ^ cw[1584] ^ cw[1586] ^ cw[1588] ^ cw[1590] ^ cw[1593] ^ cw[1595] ^ cw[1597] ^ cw[1599] ^ cw[1601] ^ cw[1603] ^ cw[1605] ^ cw[1607] ^ cw[1609] ^ cw[1611] ^ cw[1613] ^ cw[1615] ^ cw[1617] ^ cw[1619] ^ cw[1621] ^ cw[1623] ^ cw[1625] ^ cw[1627] ^ cw[1629] ^ cw[1631] ^ cw[1632] ^ cw[1634] ^ cw[1636] ^ cw[1638] ^ cw[1640] ^ cw[1642] ^ cw[1644] ^ cw[1646] ^ cw[1648] ^ cw[1650] ^ cw[1652] ^ cw[1654] ^ cw[1656] ^ cw[1658] ^ cw[1660] ^ cw[1663] ^ cw[1665] ^ cw[1667] ^ cw[1669] ^ cw[1671] ^ cw[1673] ^ cw[1675] ^ cw[1677] ^ cw[1679] ^ cw[1681] ^ cw[1683] ^ cw[1685] ^ cw[1687] ^ cw[1689] ^ cw[1691] ^ cw[1693] ^ cw[1695] ^ cw[1697] ^ cw[1699] ^ cw[1701] ^ cw[1702] ^ cw[1704] ^ cw[1706] ^ cw[1708] ^ cw[1710] ^ cw[1712] ^ cw[1714] ^ cw[1716] ^ cw[1718] ^ cw[1720] ^ cw[1722] ^ cw[1724] ^ cw[1726] ^ cw[1728] ^ cw[1730] ^ cw[1732] ^ cw[1734] ^ cw[1736] ^ cw[1738] ^ cw[1740] ^ cw[1743] ^ cw[1745] ^ cw[1747] ^ cw[1749] ^ cw[1751] ^ cw[1753] ^ cw[1755] ^ cw[1757] ^ cw[1759] ^ cw[1761] ^ cw[1763] ^ cw[1765] ^ cw[1767] ^ cw[1769] ^ cw[1771] ^ cw[1772] ^ cw[1774] ^ cw[1776] ^ cw[1778] ^ cw[1780] ^ cw[1782] ^ cw[1784] ^ cw[1786] ^ cw[1788] ^ cw[1790] ^ cw[1792] ^ cw[1794] ^ cw[1796] ^ cw[1798] ^ cw[1800] ^ cw[1803] ^ cw[1805] ^ cw[1807] ^ cw[1809] ^ cw[1811] ^ cw[1813] ^ cw[1815] ^ cw[1817] ^ cw[1819] ^ cw[1821] ^ cw[1823] ^ cw[1825] ^ cw[1827] ^ cw[1829] ^ cw[1831] ^ cw[1833] ^ cw[1835] ^ cw[1837] ^ cw[1839] ^ cw[1841] ^ cw[1842] ^ cw[1844] ^ cw[1846] ^ cw[1848] ^ cw[1850] ^ cw[1852] ^ cw[1854] ^ cw[1856] ^ cw[1858] ^ cw[1860] ^ cw[1862] ^ cw[1864] ^ cw[1866] ^ cw[1868] ^ cw[1870] ^ cw[1872] ^ cw[1874] ^ cw[1876] ^ cw[1878] ^ cw[1880] ^ cw[1883] ^ cw[1885] ^ cw[1887] ^ cw[1889] ^ cw[1891] ^ cw[1893] ^ cw[1895] ^ cw[1897] ^ cw[1899] ^ cw[1901] ^ cw[1903] ^ cw[1905] ^ cw[1907] ^ cw[1909] ^ cw[1911] ^ cw[1912] ^ cw[1914] ^ cw[1916] ^ cw[1918] ^ cw[1920] ^ cw[1922] ^ cw[1924] ^ cw[1926] ^ cw[1928] ^ cw[1930] ^ cw[1932] ^ cw[1934] ^ cw[1936] ^ cw[1938] ^ cw[1940] ^ cw[1942] ^ cw[1944] ^ cw[1946] ^ cw[1948] ^ cw[1950] ^ cw[1953] ^ cw[1955] ^ cw[1957] ^ cw[1959] ^ cw[1961] ^ cw[1963] ^ cw[1965] ^ cw[1967] ^ cw[1969] ^ cw[1971] ^ cw[1973] ^ cw[1975] ^ cw[1977] ^ cw[1979] ^ cw[1981] ^ cw[1982] ^ cw[1984] ^ cw[1986] ^ cw[1988] ^ cw[1990] ^ cw[1992] ^ cw[1994] ^ cw[1996] ^ cw[1998] ^ cw[2000] ^ cw[2002] ^ cw[2004] ^ cw[2006] ^ cw[2008] ^ cw[2010] ^ cw[2013] ^ cw[2015] ^ cw[2017] ^ cw[2019] ^ cw[2021] ^ cw[2023] ^ cw[2024] ^ cw[2025] ^ cw[2026] ^ cw[2027] ^ cw[2028] ^ cw[2029] ^ cw[2031] ^ cw[2032] ^ cw[2033] ^ cw[2034] ^ cw[2035] ^ cw[2042];
    assign syndrome[4] = cw[1] ^ cw[3] ^ cw[4] ^ cw[7] ^ cw[9] ^ cw[11] ^ cw[13] ^ cw[15] ^ cw[17] ^ cw[19] ^ cw[21] ^ cw[22] ^ cw[25] ^ cw[27] ^ cw[29] ^ cw[31] ^ cw[33] ^ cw[35] ^ cw[37] ^ cw[38] ^ cw[41] ^ cw[43] ^ cw[45] ^ cw[47] ^ cw[49] ^ cw[51] ^ cw[53] ^ cw[54] ^ cw[56] ^ cw[58] ^ cw[60] ^ cw[62] ^ cw[64] ^ cw[66] ^ cw[69] ^ cw[71] ^ cw[73] ^ cw[75] ^ cw[77] ^ cw[79] ^ cw[81] ^ cw[83] ^ cw[85] ^ cw[87] ^ cw[89] ^ cw[91] ^ cw[93] ^ cw[95] ^ cw[97] ^ cw[99] ^ cw[101] ^ cw[103] ^ cw[105] ^ cw[107] ^ cw[109] ^ cw[111] ^ cw[112] ^ cw[115] ^ cw[117] ^ cw[119] ^ cw[121] ^ cw[123] ^ cw[125] ^ cw[127] ^ cw[128] ^ cw[131] ^ cw[133] ^ cw[135] ^ cw[137] ^ cw[139] ^ cw[141] ^ cw[143] ^ cw[144] ^ cw[146] ^ cw[148] ^ cw[150] ^ cw[152] ^ cw[154] ^ cw[156] ^ cw[159] ^ cw[161] ^ cw[163] ^ cw[165] ^ cw[167] ^ cw[169] ^ cw[171] ^ cw[173] ^ cw[175] ^ cw[177] ^ cw[179] ^ cw[181] ^ cw[183] ^ cw[185] ^ cw[187] ^ cw[189] ^ cw[191] ^ cw[193] ^ cw[195] ^ cw[197] ^ cw[199] ^ cw[200] ^ cw[203] ^ cw[205] ^ cw[207] ^ cw[209] ^ cw[211] ^ cw[213] ^ cw[215] ^ cw[216] ^ cw[218] ^ cw[220] ^ cw[222] ^ cw[224] ^ cw[226] ^ cw[228] ^ cw[231] ^ cw[233] ^ cw[235] ^ cw[237] ^ cw[239] ^ cw[241] ^ cw[243] ^ cw[245] ^ cw[247] ^ cw[249] ^ cw[251] ^ cw[253] ^ cw[255] ^ cw[257] ^ cw[259] ^ cw[261] ^ cw[263] ^ cw[265] ^ cw[267] ^ cw[269] ^ cw[271] ^ cw[272] ^ cw[274] ^ cw[276] ^ cw[278] ^ cw[280] ^ cw[282] ^ cw[284] ^ cw[287] ^ cw[289] ^ cw[291] ^ cw[293] ^ cw[295] ^ cw[297] ^ cw[299] ^ cw[301] ^ cw[303] ^ cw[305] ^ cw[307] ^ cw[309] ^ cw[311] ^ cw[313] ^ cw[315] ^ cw[317] ^ cw[319] ^ cw[321] ^ cw[323] ^ cw[325] ^ cw[327] ^ cw[328] ^ cw[330] ^ cw[332] ^ cw[334] ^ cw[336] ^ cw[338] ^ cw[340] ^ cw[342] ^ cw[344] ^ cw[346] ^ cw[348] ^ cw[350] ^ cw[352] ^ cw[354] ^ cw[356] ^ cw[358] ^ cw[360] ^ cw[362] ^ cw[364] ^ cw[366] ^ cw[368] ^ cw[371] ^ cw[373] ^ cw[375] ^ cw[377] ^ cw[379] ^ cw[381] ^ cw[383] ^ cw[385] ^ cw[387] ^ cw[389] ^ cw[391] ^ cw[393] ^ cw[395] ^ cw[397] ^ cw[399] ^ cw[401] ^ cw[403] ^ cw[405] ^ cw[407] ^ cw[409] ^ cw[411] ^ cw[413] ^ cw[415] ^ cw[417] ^ cw[419] ^ cw[421] ^ cw[423] ^ cw[425] ^ cw[427] ^ cw[429] ^ cw[431] ^ cw[433] ^ cw[435] ^ cw[437] ^ cw[439] ^ cw[440] ^ cw[443] ^ cw[445] ^ cw[447] ^ cw[449] ^ cw[451] ^ cw[453] ^ cw[455] ^ cw[456] ^ cw[458] ^ cw[460] ^ cw[462] ^ cw[464] ^ cw[466] ^ cw[468] ^ cw[471] ^ cw[473] ^ cw[475] ^ cw[477] ^ cw[479] ^ cw[481] ^ cw[483] ^ cw[485] ^ cw[487] ^ cw[489] ^ cw[491] ^ cw[493] ^ cw[495] ^ cw[497] ^ cw[499] ^ cw[501] ^ cw[503] ^ cw[505] ^ cw[507] ^ cw[509] ^ cw[511] ^ cw[512] ^ cw[514] ^ cw[516] ^ cw[518] ^ cw[520] ^ cw[522] ^ cw[524] ^ cw[527] ^ cw[529] ^ cw[531] ^ cw[533] ^ cw[535] ^ cw[537] ^ cw[539] ^ cw[541] ^ cw[543] ^ cw[545] ^ cw[547] ^ cw[549] ^ cw[551] ^ cw[553] ^ cw[555] ^ cw[557] ^ cw[559] ^ cw[561] ^ cw[563] ^ cw[565] ^ cw[567] ^ cw[568] ^ cw[570] ^ cw[572] ^ cw[574] ^ cw[576] ^ cw[578] ^ cw[580] ^ cw[582] ^ cw[584] ^ cw[586] ^ cw[588] ^ cw[590] ^ cw[592] ^ cw[594] ^ cw[596] ^ cw[598] ^ cw[600] ^ cw[602] ^ cw[604] ^ cw[606] ^ cw[608] ^ cw[611] ^ cw[613] ^ cw[615] ^ cw[617] ^ cw[619] ^ cw[621] ^ cw[623] ^ cw[625] ^ cw[627] ^ cw[629] ^ cw[631] ^ cw[633] ^ cw[635] ^ cw[637] ^ cw[639] ^ cw[641] ^ cw[643] ^ cw[645] ^ cw[647] ^ cw[649] ^ cw[651] ^ cw[653] ^ cw[655] ^ cw[657] ^ cw[659] ^ cw[661] ^ cw[663] ^ cw[665] ^ cw[667] ^ cw[669] ^ cw[671] ^ cw[673] ^ cw[675] ^ cw[677] ^ cw[679] ^ cw[680] ^ cw[682] ^ cw[684] ^ cw[686] ^ cw[688] ^ cw[690] ^ cw[692] ^ cw[695] ^ cw[697] ^ cw[699] ^ cw[701] ^ cw[703] ^ cw[705] ^ cw[707] ^ cw[709] ^ cw[711] ^ cw[713] ^ cw[715] ^ cw[717] ^ cw[719] ^ cw[721] ^ cw[723] ^ cw[725] ^ cw[727] ^ cw[729] ^ cw[731] ^ cw[733] ^ cw[735] ^ cw[736] ^ cw[738] ^ cw[740] ^ cw[742] ^ cw[744] ^ cw[746] ^ cw[748] ^ cw[750] ^ cw[752] ^ cw[754] ^ cw[756] ^ cw[758] ^ cw[760] ^ cw[762] ^ cw[764] ^ cw[766] ^ cw[768] ^ cw[770] ^ cw[772] ^ cw[774] ^ cw[776] ^ cw[779] ^ cw[781] ^ cw[783] ^ cw[785] ^ cw[787] ^ cw[789] ^ cw[791] ^ cw[793] ^ cw[795] ^ cw[797] ^ cw[799] ^ cw[801] ^ cw[803] ^ cw[805] ^ cw[807] ^ cw[809] ^ cw[811] ^ cw[813] ^ cw[815] ^ cw[817] ^ cw[819] ^ cw[821] ^ cw[823] ^ cw[825] ^ cw[827] ^ cw[829] ^ cw[831] ^ cw[833] ^ cw[835] ^ cw[837] ^ cw[839] ^ cw[841] ^ cw[843] ^ cw[845] ^ cw[847] ^ cw[848] ^ cw[850] ^ cw[852] ^ cw[854] ^ cw[856] ^ cw[858] ^ cw[860] ^ cw[862] ^ cw[864] ^ cw[866] ^ cw[868] ^ cw[870] ^ cw[872] ^ cw[874] ^ cw[876] ^ cw[878] ^ cw[880] ^ cw[882] ^ cw[884] ^ cw[886] ^ cw[888] ^ cw[891] ^ cw[893] ^ cw[895] ^ cw[897] ^ cw[899] ^ cw[901] ^ cw[903] ^ cw[905] ^ cw[907] ^ cw[909] ^ cw[911] ^ cw[913] ^ cw[915] ^ cw[917] ^ cw[919] ^ cw[921] ^ cw[923] ^ cw[925] ^ cw[927] ^ cw[929] ^ cw[931] ^ cw[933] ^ cw[935] ^ cw[937] ^ cw[939] ^ cw[941] ^ cw[943] ^ cw[945] ^ cw[947] ^ cw[949] ^ cw[951] ^ cw[953] ^ cw[955] ^ cw[957] ^ cw[959] ^ cw[960] ^ cw[962] ^ cw[964] ^ cw[966] ^ cw[968] ^ cw[970] ^ cw[972] ^ cw[974] ^ cw[976] ^ cw[978] ^ cw[980] ^ cw[982] ^ cw[984] ^ cw[986] ^ cw[988] ^ cw[990] ^ cw[992] ^ cw[994] ^ cw[996] ^ cw[998] ^ cw[1000] ^ cw[1002] ^ cw[1004] ^ cw[1006] ^ cw[1008] ^ cw[1010] ^ cw[1012] ^ cw[1014] ^ cw[1016] ^ cw[1018] ^ cw[1020] ^ cw[1022] ^ cw[1024] ^ cw[1026] ^ cw[1028] ^ cw[1031] ^ cw[1033] ^ cw[1035] ^ cw[1037] ^ cw[1039] ^ cw[1041] ^ cw[1043] ^ cw[1045] ^ cw[1047] ^ cw[1049] ^ cw[1051] ^ cw[1053] ^ cw[1055] ^ cw[1057] ^ cw[1059] ^ cw[1061] ^ cw[1063] ^ cw[1065] ^ cw[1067] ^ cw[1069] ^ cw[1071] ^ cw[1073] ^ cw[1075] ^ cw[1077] ^ cw[1079] ^ cw[1081] ^ cw[1083] ^ cw[1085] ^ cw[1087] ^ cw[1089] ^ cw[1091] ^ cw[1093] ^ cw[1095] ^ cw[1097] ^ cw[1099] ^ cw[1100] ^ cw[1102] ^ cw[1104] ^ cw[1106] ^ cw[1108] ^ cw[1110] ^ cw[1112] ^ cw[1115] ^ cw[1117] ^ cw[1119] ^ cw[1121] ^ cw[1123] ^ cw[1125] ^ cw[1127] ^ cw[1129] ^ cw[1131] ^ cw[1133] ^ cw[1135] ^ cw[1137] ^ cw[1139] ^ cw[1141] ^ cw[1143] ^ cw[1145] ^ cw[1147] ^ cw[1149] ^ cw[1151] ^ cw[1153] ^ cw[1155] ^ cw[1156] ^ cw[1158] ^ cw[1160] ^ cw[1162] ^ cw[1164] ^ cw[1166] ^ cw[1168] ^ cw[1170] ^ cw[1172] ^ cw[1174] ^ cw[1176] ^ cw[1178] ^ cw[1180] ^ cw[1182] ^ cw[1184] ^ cw[1186] ^ cw[1188] ^ cw[1190] ^ cw[1192] ^ cw[1194] ^ cw[1196] ^ cw[1199] ^ cw[1201] ^ cw[1203] ^ cw[1205] ^ cw[1207] ^ cw[1209] ^ cw[1211] ^ cw[1213] ^ cw[1215] ^ cw[1217] ^ cw[1219] ^ cw[1221] ^ cw[1223] ^ cw[1225] ^ cw[1227] ^ cw[1229] ^ cw[1231] ^ cw[1233] ^ cw[1235] ^ cw[1237] ^ cw[1239] ^ cw[1241] ^ cw[1243] ^ cw[1245] ^ cw[1247] ^ cw[1249] ^ cw[1251] ^ cw[1253] ^ cw[1255] ^ cw[1257] ^ cw[1259] ^ cw[1261] ^ cw[1263] ^ cw[1265] ^ cw[1267] ^ cw[1268] ^ cw[1270] ^ cw[1272] ^ cw[1274] ^ cw[1276] ^ cw[1278] ^ cw[1280] ^ cw[1282] ^ cw[1284] ^ cw[1286] ^ cw[1288] ^ cw[1290] ^ cw[1292] ^ cw[1294] ^ cw[1296] ^ cw[1298] ^ cw[1300] ^ cw[1302] ^ cw[1304] ^ cw[1306] ^ cw[1308] ^ cw[1311] ^ cw[1313] ^ cw[1315] ^ cw[1317] ^ cw[1319] ^ cw[1321] ^ cw[1323] ^ cw[1325] ^ cw[1327] ^ cw[1329] ^ cw[1331] ^ cw[1333] ^ cw[1335] ^ cw[1337] ^ cw[1339] ^ cw[1341] ^ cw[1343] ^ cw[1345] ^ cw[1347] ^ cw[1349] ^ cw[1351] ^ cw[1353] ^ cw[1355] ^ cw[1357] ^ cw[1359] ^ cw[1361] ^ cw[1363] ^ cw[1365] ^ cw[1367] ^ cw[1369] ^ cw[1371] ^ cw[1373] ^ cw[1375] ^ cw[1377] ^ cw[1379] ^ cw[1380] ^ cw[1382] ^ cw[1384] ^ cw[1386] ^ cw[1388] ^ cw[1390] ^ cw[1392] ^ cw[1394] ^ cw[1396] ^ cw[1398] ^ cw[1400] ^ cw[1402] ^ cw[1404] ^ cw[1406] ^ cw[1408] ^ cw[1410] ^ cw[1412] ^ cw[1414] ^ cw[1416] ^ cw[1418] ^ cw[1420] ^ cw[1422] ^ cw[1424] ^ cw[1426] ^ cw[1428] ^ cw[1430] ^ cw[1432] ^ cw[1434] ^ cw[1436] ^ cw[1438] ^ cw[1440] ^ cw[1442] ^ cw[1444] ^ cw[1446] ^ cw[1448] ^ cw[1451] ^ cw[1453] ^ cw[1455] ^ cw[1457] ^ cw[1459] ^ cw[1461] ^ cw[1463] ^ cw[1465] ^ cw[1467] ^ cw[1469] ^ cw[1471] ^ cw[1473] ^ cw[1475] ^ cw[1477] ^ cw[1479] ^ cw[1481] ^ cw[1483] ^ cw[1485] ^ cw[1487] ^ cw[1489] ^ cw[1491] ^ cw[1493] ^ cw[1495] ^ cw[1497] ^ cw[1499] ^ cw[1501] ^ cw[1503] ^ cw[1505] ^ cw[1507] ^ cw[1509] ^ cw[1511] ^ cw[1513] ^ cw[1515] ^ cw[1517] ^ cw[1519] ^ cw[1520] ^ cw[1522] ^ cw[1524] ^ cw[1526] ^ cw[1528] ^ cw[1530] ^ cw[1532] ^ cw[1534] ^ cw[1536] ^ cw[1538] ^ cw[1540] ^ cw[1542] ^ cw[1544] ^ cw[1546] ^ cw[1548] ^ cw[1550] ^ cw[1552] ^ cw[1554] ^ cw[1556] ^ cw[1558] ^ cw[1560] ^ cw[1563] ^ cw[1565] ^ cw[1567] ^ cw[1569] ^ cw[1571] ^ cw[1573] ^ cw[1575] ^ cw[1577] ^ cw[1579] ^ cw[1581] ^ cw[1583] ^ cw[1585] ^ cw[1587] ^ cw[1589] ^ cw[1591] ^ cw[1593] ^ cw[1595] ^ cw[1597] ^ cw[1599] ^ cw[1601] ^ cw[1603] ^ cw[1605] ^ cw[1607] ^ cw[1609] ^ cw[1611] ^ cw[1613] ^ cw[1615] ^ cw[1617] ^ cw[1619] ^ cw[1621] ^ cw[1623] ^ cw[1625] ^ cw[1627] ^ cw[1629] ^ cw[1631] ^ cw[1632] ^ cw[1634] ^ cw[1636] ^ cw[1638] ^ cw[1640] ^ cw[1642] ^ cw[1644] ^ cw[1646] ^ cw[1648] ^ cw[1650] ^ cw[1652] ^ cw[1654] ^ cw[1656] ^ cw[1658] ^ cw[1660] ^ cw[1662] ^ cw[1664] ^ cw[1666] ^ cw[1668] ^ cw[1670] ^ cw[1672] ^ cw[1674] ^ cw[1676] ^ cw[1678] ^ cw[1680] ^ cw[1682] ^ cw[1684] ^ cw[1686] ^ cw[1688] ^ cw[1690] ^ cw[1692] ^ cw[1694] ^ cw[1696] ^ cw[1698] ^ cw[1700] ^ cw[1703] ^ cw[1705] ^ cw[1707] ^ cw[1709] ^ cw[1711] ^ cw[1713] ^ cw[1715] ^ cw[1717] ^ cw[1719] ^ cw[1721] ^ cw[1723] ^ cw[1725] ^ cw[1727] ^ cw[1729] ^ cw[1731] ^ cw[1733] ^ cw[1735] ^ cw[1737] ^ cw[1739] ^ cw[1741] ^ cw[1743] ^ cw[1745] ^ cw[1747] ^ cw[1749] ^ cw[1751] ^ cw[1753] ^ cw[1755] ^ cw[1757] ^ cw[1759] ^ cw[1761] ^ cw[1763] ^ cw[1765] ^ cw[1767] ^ cw[1769] ^ cw[1771] ^ cw[1772] ^ cw[1774] ^ cw[1776] ^ cw[1778] ^ cw[1780] ^ cw[1782] ^ cw[1784] ^ cw[1786] ^ cw[1788] ^ cw[1790] ^ cw[1792] ^ cw[1794] ^ cw[1796] ^ cw[1798] ^ cw[1800] ^ cw[1802] ^ cw[1804] ^ cw[1806] ^ cw[1808] ^ cw[1810] ^ cw[1812] ^ cw[1814] ^ cw[1816] ^ cw[1818] ^ cw[1820] ^ cw[1822] ^ cw[1824] ^ cw[1826] ^ cw[1828] ^ cw[1830] ^ cw[1832] ^ cw[1834] ^ cw[1836] ^ cw[1838] ^ cw[1840] ^ cw[1843] ^ cw[1845] ^ cw[1847] ^ cw[1849] ^ cw[1851] ^ cw[1853] ^ cw[1855] ^ cw[1857] ^ cw[1859] ^ cw[1861] ^ cw[1863] ^ cw[1865] ^ cw[1867] ^ cw[1869] ^ cw[1871] ^ cw[1873] ^ cw[1875] ^ cw[1877] ^ cw[1879] ^ cw[1881] ^ cw[1883] ^ cw[1885] ^ cw[1887] ^ cw[1889] ^ cw[1891] ^ cw[1893] ^ cw[1895] ^ cw[1897] ^ cw[1899] ^ cw[1901] ^ cw[1903] ^ cw[1905] ^ cw[1907] ^ cw[1909] ^ cw[1911] ^ cw[1912] ^ cw[1914] ^ cw[1916] ^ cw[1918] ^ cw[1920] ^ cw[1922] ^ cw[1924] ^ cw[1926] ^ cw[1928] ^ cw[1930] ^ cw[1932] ^ cw[1934] ^ cw[1936] ^ cw[1938] ^ cw[1940] ^ cw[1942] ^ cw[1944] ^ cw[1946] ^ cw[1948] ^ cw[1950] ^ cw[1952] ^ cw[1954] ^ cw[1956] ^ cw[1958] ^ cw[1960] ^ cw[1962] ^ cw[1964] ^ cw[1966] ^ cw[1968] ^ cw[1970] ^ cw[1972] ^ cw[1974] ^ cw[1976] ^ cw[1978] ^ cw[1980] ^ cw[1983] ^ cw[1985] ^ cw[1987] ^ cw[1989] ^ cw[1991] ^ cw[1993] ^ cw[1995] ^ cw[1997] ^ cw[1999] ^ cw[2001] ^ cw[2003] ^ cw[2005] ^ cw[2007] ^ cw[2009] ^ cw[2011] ^ cw[2013] ^ cw[2015] ^ cw[2017] ^ cw[2019] ^ cw[2021] ^ cw[2023] ^ cw[2024] ^ cw[2025] ^ cw[2026] ^ cw[2027] ^ cw[2028] ^ cw[2029] ^ cw[2030] ^ cw[2032] ^ cw[2033] ^ cw[2034] ^ cw[2035] ^ cw[2043];
    assign syndrome[3] = cw[1] ^ cw[2] ^ cw[5] ^ cw[7] ^ cw[9] ^ cw[11] ^ cw[13] ^ cw[15] ^ cw[17] ^ cw[19] ^ cw[20] ^ cw[23] ^ cw[25] ^ cw[27] ^ cw[29] ^ cw[31] ^ cw[33] ^ cw[35] ^ cw[37] ^ cw[38] ^ cw[40] ^ cw[42] ^ cw[44] ^ cw[46] ^ cw[48] ^ cw[50] ^ cw[52] ^ cw[55] ^ cw[57] ^ cw[59] ^ cw[61] ^ cw[63] ^ cw[65] ^ cw[67] ^ cw[69] ^ cw[71] ^ cw[73] ^ cw[75] ^ cw[77] ^ cw[79] ^ cw[81] ^ cw[83] ^ cw[85] ^ cw[87] ^ cw[89] ^ cw[91] ^ cw[93] ^ cw[95] ^ cw[97] ^ cw[99] ^ cw[101] ^ cw[103] ^ cw[105] ^ cw[107] ^ cw[109] ^ cw[110] ^ cw[113] ^ cw[115] ^ cw[117] ^ cw[119] ^ cw[121] ^ cw[123] ^ cw[125] ^ cw[127] ^ cw[128] ^ cw[130] ^ cw[132] ^ cw[134] ^ cw[136] ^ cw[138] ^ cw[140] ^ cw[142] ^ cw[145] ^ cw[147] ^ cw[149] ^ cw[151] ^ cw[153] ^ cw[155] ^ cw[157] ^ cw[159] ^ cw[161] ^ cw[163] ^ cw[165] ^ cw[167] ^ cw[169] ^ cw[171] ^ cw[173] ^ cw[175] ^ cw[177] ^ cw[179] ^ cw[181] ^ cw[183] ^ cw[185] ^ cw[187] ^ cw[189] ^ cw[191] ^ cw[193] ^ cw[195] ^ cw[197] ^ cw[199] ^ cw[200] ^ cw[202] ^ cw[204] ^ cw[206] ^ cw[208] ^ cw[210] ^ cw[212] ^ cw[214] ^ cw[217] ^ cw[219] ^ cw[221] ^ cw[223] ^ cw[225] ^ cw[227] ^ cw[229] ^ cw[231] ^ cw[233] ^ cw[235] ^ cw[237] ^ cw[239] ^ cw[241] ^ cw[243] ^ cw[245] ^ cw[247] ^ cw[249] ^ cw[251] ^ cw[253] ^ cw[255] ^ cw[257] ^ cw[259] ^ cw[261] ^ cw[263] ^ cw[265] ^ cw[267] ^ cw[269] ^ cw[271] ^ cw[272] ^ cw[274] ^ cw[276] ^ cw[278] ^ cw[280] ^ cw[282] ^ cw[284] ^ cw[286] ^ cw[288] ^ cw[290] ^ cw[292] ^ cw[294] ^ cw[296] ^ cw[298] ^ cw[300] ^ cw[302] ^ cw[304] ^ cw[306] ^ cw[308] ^ cw[310] ^ cw[312] ^ cw[314] ^ cw[316] ^ cw[318] ^ cw[320] ^ cw[322] ^ cw[324] ^ cw[326] ^ cw[329] ^ cw[331] ^ cw[333] ^ cw[335] ^ cw[337] ^ cw[339] ^ cw[341] ^ cw[343] ^ cw[345] ^ cw[347] ^ cw[349] ^ cw[351] ^ cw[353] ^ cw[355] ^ cw[357] ^ cw[359] ^ cw[361] ^ cw[363] ^ cw[365] ^ cw[367] ^ cw[369] ^ cw[371] ^ cw[373] ^ cw[375] ^ cw[377] ^ cw[379] ^ cw[381] ^ cw[383] ^ cw[385] ^ cw[387] ^ cw[389] ^ cw[391] ^ cw[393] ^ cw[395] ^ cw[397] ^ cw[399] ^ cw[401] ^ cw[403] ^ cw[405] ^ cw[407] ^ cw[409] ^ cw[411] ^ cw[413] ^ cw[415] ^ cw[417] ^ cw[419] ^ cw[421] ^ cw[423] ^ cw[425] ^ cw[427] ^ cw[429] ^ cw[431] ^ cw[433] ^ cw[435] ^ cw[437] ^ cw[439] ^ cw[440] ^ cw[442] ^ cw[444] ^ cw[446] ^ cw[448] ^ cw[450] ^ cw[452] ^ cw[454] ^ cw[457] ^ cw[459] ^ cw[461] ^ cw[463] ^ cw[465] ^ cw[467] ^ cw[469] ^ cw[471] ^ cw[473] ^ cw[475] ^ cw[477] ^ cw[479] ^ cw[481] ^ cw[483] ^ cw[485] ^ cw[487] ^ cw[489] ^ cw[491] ^ cw[493] ^ cw[495] ^ cw[497] ^ cw[499] ^ cw[501] ^ cw[503] ^ cw[505] ^ cw[507] ^ cw[509] ^ cw[511] ^ cw[512] ^ cw[514] ^ cw[516] ^ cw[518] ^ cw[520] ^ cw[522] ^ cw[524] ^ cw[526] ^ cw[528] ^ cw[530] ^ cw[532] ^ cw[534] ^ cw[536] ^ cw[538] ^ cw[540] ^ cw[542] ^ cw[544] ^ cw[546] ^ cw[548] ^ cw[550] ^ cw[552] ^ cw[554] ^ cw[556] ^ cw[558] ^ cw[560] ^ cw[562] ^ cw[564] ^ cw[566] ^ cw[569] ^ cw[571] ^ cw[573] ^ cw[575] ^ cw[577] ^ cw[579] ^ cw[581] ^ cw[583] ^ cw[585] ^ cw[587] ^ cw[589] ^ cw[591] ^ cw[593] ^ cw[595] ^ cw[597] ^ cw[599] ^ cw[601] ^ cw[603] ^ cw[605] ^ cw[607] ^ cw[609] ^ cw[611] ^ cw[613] ^ cw[615] ^ cw[617] ^ cw[619] ^ cw[621] ^ cw[623] ^ cw[625] ^ cw[627] ^ cw[629] ^ cw[631] ^ cw[633] ^ cw[635] ^ cw[637] ^ cw[639] ^ cw[641] ^ cw[643] ^ cw[645] ^ cw[647] ^ cw[649] ^ cw[651] ^ cw[653] ^ cw[655] ^ cw[657] ^ cw[659] ^ cw[661] ^ cw[663] ^ cw[665] ^ cw[667] ^ cw[669] ^ cw[671] ^ cw[673] ^ cw[675] ^ cw[677] ^ cw[679] ^ cw[680] ^ cw[682] ^ cw[684] ^ cw[686] ^ cw[688] ^ cw[690] ^ cw[692] ^ cw[694] ^ cw[696] ^ cw[698] ^ cw[700] ^ cw[702] ^ cw[704] ^ cw[706] ^ cw[708] ^ cw[710] ^ cw[712] ^ cw[714] ^ cw[716] ^ cw[718] ^ cw[720] ^ cw[722] ^ cw[724] ^ cw[726] ^ cw[728] ^ cw[730] ^ cw[732] ^ cw[734] ^ cw[737] ^ cw[739] ^ cw[741] ^ cw[743] ^ cw[745] ^ cw[747] ^ cw[749] ^ cw[751] ^ cw[753] ^ cw[755] ^ cw[757] ^ cw[759] ^ cw[761] ^ cw[763] ^ cw[765] ^ cw[767] ^ cw[769] ^ cw[771] ^ cw[773] ^ cw[775] ^ cw[777] ^ cw[779] ^ cw[781] ^ cw[783] ^ cw[785] ^ cw[787] ^ cw[789] ^ cw[791] ^ cw[793] ^ cw[795] ^ cw[797] ^ cw[799] ^ cw[801] ^ cw[803] ^ cw[805] ^ cw[807] ^ cw[809] ^ cw[811] ^ cw[813] ^ cw[815] ^ cw[817] ^ cw[819] ^ cw[821] ^ cw[823] ^ cw[825] ^ cw[827] ^ cw[829] ^ cw[831] ^ cw[833] ^ cw[835] ^ cw[837] ^ cw[839] ^ cw[841] ^ cw[843] ^ cw[845] ^ cw[847] ^ cw[848] ^ cw[850] ^ cw[852] ^ cw[854] ^ cw[856] ^ cw[858] ^ cw[860] ^ cw[862] ^ cw[864] ^ cw[866] ^ cw[868] ^ cw[870] ^ cw[872] ^ cw[874] ^ cw[876] ^ cw[878] ^ cw[880] ^ cw[882] ^ cw[884] ^ cw[886] ^ cw[888] ^ cw[890] ^ cw[892] ^ cw[894] ^ cw[896] ^ cw[898] ^ cw[900] ^ cw[902] ^ cw[904] ^ cw[906] ^ cw[908] ^ cw[910] ^ cw[912] ^ cw[914] ^ cw[916] ^ cw[918] ^ cw[920] ^ cw[922] ^ cw[924] ^ cw[926] ^ cw[928] ^ cw[930] ^ cw[932] ^ cw[934] ^ cw[936] ^ cw[938] ^ cw[940] ^ cw[942] ^ cw[944] ^ cw[946] ^ cw[948] ^ cw[950] ^ cw[952] ^ cw[954] ^ cw[956] ^ cw[958] ^ cw[961] ^ cw[963] ^ cw[965] ^ cw[967] ^ cw[969] ^ cw[971] ^ cw[973] ^ cw[975] ^ cw[977] ^ cw[979] ^ cw[981] ^ cw[983] ^ cw[985] ^ cw[987] ^ cw[989] ^ cw[991] ^ cw[993] ^ cw[995] ^ cw[997] ^ cw[999] ^ cw[1001] ^ cw[1003] ^ cw[1005] ^ cw[1007] ^ cw[1009] ^ cw[1011] ^ cw[1013] ^ cw[1015] ^ cw[1017] ^ cw[1019] ^ cw[1021] ^ cw[1023] ^ cw[1025] ^ cw[1027] ^ cw[1029] ^ cw[1031] ^ cw[1033] ^ cw[1035] ^ cw[1037] ^ cw[1039] ^ cw[1041] ^ cw[1043] ^ cw[1045] ^ cw[1047] ^ cw[1049] ^ cw[1051] ^ cw[1053] ^ cw[1055] ^ cw[1057] ^ cw[1059] ^ cw[1061] ^ cw[1063] ^ cw[1065] ^ cw[1067] ^ cw[1069] ^ cw[1071] ^ cw[1073] ^ cw[1075] ^ cw[1077] ^ cw[1079] ^ cw[1081] ^ cw[1083] ^ cw[1085] ^ cw[1087] ^ cw[1089] ^ cw[1091] ^ cw[1093] ^ cw[1095] ^ cw[1097] ^ cw[1099] ^ cw[1100] ^ cw[1102] ^ cw[1104] ^ cw[1106] ^ cw[1108] ^ cw[1110] ^ cw[1112] ^ cw[1114] ^ cw[1116] ^ cw[1118] ^ cw[1120] ^ cw[1122] ^ cw[1124] ^ cw[1126] ^ cw[1128] ^ cw[1130] ^ cw[1132] ^ cw[1134] ^ cw[1136] ^ cw[1138] ^ cw[1140] ^ cw[1142] ^ cw[1144] ^ cw[1146] ^ cw[1148] ^ cw[1150] ^ cw[1152] ^ cw[1154] ^ cw[1157] ^ cw[1159] ^ cw[1161] ^ cw[1163] ^ cw[1165] ^ cw[1167] ^ cw[1169] ^ cw[1171] ^ cw[1173] ^ cw[1175] ^ cw[1177] ^ cw[1179] ^ cw[1181] ^ cw[1183] ^ cw[1185] ^ cw[1187] ^ cw[1189] ^ cw[1191] ^ cw[1193] ^ cw[1195] ^ cw[1197] ^ cw[1199] ^ cw[1201] ^ cw[1203] ^ cw[1205] ^ cw[1207] ^ cw[1209] ^ cw[1211] ^ cw[1213] ^ cw[1215] ^ cw[1217] ^ cw[1219] ^ cw[1221] ^ cw[1223] ^ cw[1225] ^ cw[1227] ^ cw[1229] ^ cw[1231] ^ cw[1233] ^ cw[1235] ^ cw[1237] ^ cw[1239] ^ cw[1241] ^ cw[1243] ^ cw[1245] ^ cw[1247] ^ cw[1249] ^ cw[1251] ^ cw[1253] ^ cw[1255] ^ cw[1257] ^ cw[1259] ^ cw[1261] ^ cw[1263] ^ cw[1265] ^ cw[1267] ^ cw[1268] ^ cw[1270] ^ cw[1272] ^ cw[1274] ^ cw[1276] ^ cw[1278] ^ cw[1280] ^ cw[1282] ^ cw[1284] ^ cw[1286] ^ cw[1288] ^ cw[1290] ^ cw[1292] ^ cw[1294] ^ cw[1296] ^ cw[1298] ^ cw[1300] ^ cw[1302] ^ cw[1304] ^ cw[1306] ^ cw[1308] ^ cw[1310] ^ cw[1312] ^ cw[1314] ^ cw[1316] ^ cw[1318] ^ cw[1320] ^ cw[1322] ^ cw[1324] ^ cw[1326] ^ cw[1328] ^ cw[1330] ^ cw[1332] ^ cw[1334] ^ cw[1336] ^ cw[1338] ^ cw[1340] ^ cw[1342] ^ cw[1344] ^ cw[1346] ^ cw[1348] ^ cw[1350] ^ cw[1352] ^ cw[1354] ^ cw[1356] ^ cw[1358] ^ cw[1360] ^ cw[1362] ^ cw[1364] ^ cw[1366] ^ cw[1368] ^ cw[1370] ^ cw[1372] ^ cw[1374] ^ cw[1376] ^ cw[1378] ^ cw[1381] ^ cw[1383] ^ cw[1385] ^ cw[1387] ^ cw[1389] ^ cw[1391] ^ cw[1393] ^ cw[1395] ^ cw[1397] ^ cw[1399] ^ cw[1401] ^ cw[1403] ^ cw[1405] ^ cw[1407] ^ cw[1409] ^ cw[1411] ^ cw[1413] ^ cw[1415] ^ cw[1417] ^ cw[1419] ^ cw[1421] ^ cw[1423] ^ cw[1425] ^ cw[1427] ^ cw[1429] ^ cw[1431] ^ cw[1433] ^ cw[1435] ^ cw[1437] ^ cw[1439] ^ cw[1441] ^ cw[1443] ^ cw[1445] ^ cw[1447] ^ cw[1449] ^ cw[1451] ^ cw[1453] ^ cw[1455] ^ cw[1457] ^ cw[1459] ^ cw[1461] ^ cw[1463] ^ cw[1465] ^ cw[1467] ^ cw[1469] ^ cw[1471] ^ cw[1473] ^ cw[1475] ^ cw[1477] ^ cw[1479] ^ cw[1481] ^ cw[1483] ^ cw[1485] ^ cw[1487] ^ cw[1489] ^ cw[1491] ^ cw[1493] ^ cw[1495] ^ cw[1497] ^ cw[1499] ^ cw[1501] ^ cw[1503] ^ cw[1505] ^ cw[1507] ^ cw[1509] ^ cw[1511] ^ cw[1513] ^ cw[1515] ^ cw[1517] ^ cw[1519] ^ cw[1520] ^ cw[1522] ^ cw[1524] ^ cw[1526] ^ cw[1528] ^ cw[1530] ^ cw[1532] ^ cw[1534] ^ cw[1536] ^ cw[1538] ^ cw[1540] ^ cw[1542] ^ cw[1544] ^ cw[1546] ^ cw[1548] ^ cw[1550] ^ cw[1552] ^ cw[1554] ^ cw[1556] ^ cw[1558] ^ cw[1560] ^ cw[1562] ^ cw[1564] ^ cw[1566] ^ cw[1568] ^ cw[1570] ^ cw[1572] ^ cw[1574] ^ cw[1576] ^ cw[1578] ^ cw[1580] ^ cw[1582] ^ cw[1584] ^ cw[1586] ^ cw[1588] ^ cw[1590] ^ cw[1592] ^ cw[1594] ^ cw[1596] ^ cw[1598] ^ cw[1600] ^ cw[1602] ^ cw[1604] ^ cw[1606] ^ cw[1608] ^ cw[1610] ^ cw[1612] ^ cw[1614] ^ cw[1616] ^ cw[1618] ^ cw[1620] ^ cw[1622] ^ cw[1624] ^ cw[1626] ^ cw[1628] ^ cw[1630] ^ cw[1633] ^ cw[1635] ^ cw[1637] ^ cw[1639] ^ cw[1641] ^ cw[1643] ^ cw[1645] ^ cw[1647] ^ cw[1649] ^ cw[1651] ^ cw[1653] ^ cw[1655] ^ cw[1657] ^ cw[1659] ^ cw[1661] ^ cw[1663] ^ cw[1665] ^ cw[1667] ^ cw[1669] ^ cw[1671] ^ cw[1673] ^ cw[1675] ^ cw[1677] ^ cw[1679] ^ cw[1681] ^ cw[1683] ^ cw[1685] ^ cw[1687] ^ cw[1689] ^ cw[1691] ^ cw[1693] ^ cw[1695] ^ cw[1697] ^ cw[1699] ^ cw[1701] ^ cw[1703] ^ cw[1705] ^ cw[1707] ^ cw[1709] ^ cw[1711] ^ cw[1713] ^ cw[1715] ^ cw[1717] ^ cw[1719] ^ cw[1721] ^ cw[1723] ^ cw[1725] ^ cw[1727] ^ cw[1729] ^ cw[1731] ^ cw[1733] ^ cw[1735] ^ cw[1737] ^ cw[1739] ^ cw[1741] ^ cw[1743] ^ cw[1745] ^ cw[1747] ^ cw[1749] ^ cw[1751] ^ cw[1753] ^ cw[1755] ^ cw[1757] ^ cw[1759] ^ cw[1761] ^ cw[1763] ^ cw[1765] ^ cw[1767] ^ cw[1769] ^ cw[1771] ^ cw[1772] ^ cw[1774] ^ cw[1776] ^ cw[1778] ^ cw[1780] ^ cw[1782] ^ cw[1784] ^ cw[1786] ^ cw[1788] ^ cw[1790] ^ cw[1792] ^ cw[1794] ^ cw[1796] ^ cw[1798] ^ cw[1800] ^ cw[1802] ^ cw[1804] ^ cw[1806] ^ cw[1808] ^ cw[1810] ^ cw[1812] ^ cw[1814] ^ cw[1816] ^ cw[1818] ^ cw[1820] ^ cw[1822] ^ cw[1824] ^ cw[1826] ^ cw[1828] ^ cw[1830] ^ cw[1832] ^ cw[1834] ^ cw[1836] ^ cw[1838] ^ cw[1840] ^ cw[1842] ^ cw[1844] ^ cw[1846] ^ cw[1848] ^ cw[1850] ^ cw[1852] ^ cw[1854] ^ cw[1856] ^ cw[1858] ^ cw[1860] ^ cw[1862] ^ cw[1864] ^ cw[1866] ^ cw[1868] ^ cw[1870] ^ cw[1872] ^ cw[1874] ^ cw[1876] ^ cw[1878] ^ cw[1880] ^ cw[1882] ^ cw[1884] ^ cw[1886] ^ cw[1888] ^ cw[1890] ^ cw[1892] ^ cw[1894] ^ cw[1896] ^ cw[1898] ^ cw[1900] ^ cw[1902] ^ cw[1904] ^ cw[1906] ^ cw[1908] ^ cw[1910] ^ cw[1913] ^ cw[1915] ^ cw[1917] ^ cw[1919] ^ cw[1921] ^ cw[1923] ^ cw[1925] ^ cw[1927] ^ cw[1929] ^ cw[1931] ^ cw[1933] ^ cw[1935] ^ cw[1937] ^ cw[1939] ^ cw[1941] ^ cw[1943] ^ cw[1945] ^ cw[1947] ^ cw[1949] ^ cw[1951] ^ cw[1953] ^ cw[1955] ^ cw[1957] ^ cw[1959] ^ cw[1961] ^ cw[1963] ^ cw[1965] ^ cw[1967] ^ cw[1969] ^ cw[1971] ^ cw[1973] ^ cw[1975] ^ cw[1977] ^ cw[1979] ^ cw[1981] ^ cw[1983] ^ cw[1985] ^ cw[1987] ^ cw[1989] ^ cw[1991] ^ cw[1993] ^ cw[1995] ^ cw[1997] ^ cw[1999] ^ cw[2001] ^ cw[2003] ^ cw[2005] ^ cw[2007] ^ cw[2009] ^ cw[2011] ^ cw[2013] ^ cw[2015] ^ cw[2017] ^ cw[2019] ^ cw[2021] ^ cw[2023] ^ cw[2024] ^ cw[2025] ^ cw[2026] ^ cw[2027] ^ cw[2028] ^ cw[2029] ^ cw[2030] ^ cw[2031] ^ cw[2033] ^ cw[2034] ^ cw[2035] ^ cw[2044];
    assign syndrome[2] = cw[0] ^ cw[3] ^ cw[5] ^ cw[7] ^ cw[9] ^ cw[11] ^ cw[13] ^ cw[15] ^ cw[17] ^ cw[19] ^ cw[20] ^ cw[22] ^ cw[24] ^ cw[26] ^ cw[28] ^ cw[30] ^ cw[32] ^ cw[34] ^ cw[36] ^ cw[39] ^ cw[41] ^ cw[43] ^ cw[45] ^ cw[47] ^ cw[49] ^ cw[51] ^ cw[53] ^ cw[55] ^ cw[57] ^ cw[59] ^ cw[61] ^ cw[63] ^ cw[65] ^ cw[67] ^ cw[69] ^ cw[71] ^ cw[73] ^ cw[75] ^ cw[77] ^ cw[79] ^ cw[81] ^ cw[83] ^ cw[85] ^ cw[87] ^ cw[89] ^ cw[91] ^ cw[93] ^ cw[95] ^ cw[97] ^ cw[99] ^ cw[101] ^ cw[103] ^ cw[105] ^ cw[107] ^ cw[109] ^ cw[110] ^ cw[112] ^ cw[114] ^ cw[116] ^ cw[118] ^ cw[120] ^ cw[122] ^ cw[124] ^ cw[126] ^ cw[129] ^ cw[131] ^ cw[133] ^ cw[135] ^ cw[137] ^ cw[139] ^ cw[141] ^ cw[143] ^ cw[145] ^ cw[147] ^ cw[149] ^ cw[151] ^ cw[153] ^ cw[155] ^ cw[157] ^ cw[159] ^ cw[161] ^ cw[163] ^ cw[165] ^ cw[167] ^ cw[169] ^ cw[171] ^ cw[173] ^ cw[175] ^ cw[177] ^ cw[179] ^ cw[181] ^ cw[183] ^ cw[185] ^ cw[187] ^ cw[189] ^ cw[191] ^ cw[193] ^ cw[195] ^ cw[197] ^ cw[199] ^ cw[200] ^ cw[202] ^ cw[204] ^ cw[206] ^ cw[208] ^ cw[210] ^ cw[212] ^ cw[214] ^ cw[216] ^ cw[218] ^ cw[220] ^ cw[222] ^ cw[224] ^ cw[226] ^ cw[228] ^ cw[230] ^ cw[232] ^ cw[234] ^ cw[236] ^ cw[238] ^ cw[240] ^ cw[242] ^ cw[244] ^ cw[246] ^ cw[248] ^ cw[250] ^ cw[252] ^ cw[254] ^ cw[256] ^ cw[258] ^ cw[260] ^ cw[262] ^ cw[264] ^ cw[266] ^ cw[268] ^ cw[270] ^ cw[273] ^ cw[275] ^ cw[277] ^ cw[279] ^ cw[281] ^ cw[283] ^ cw[285] ^ cw[287] ^ cw[289] ^ cw[291] ^ cw[293] ^ cw[295] ^ cw[297] ^ cw[299] ^ cw[301] ^ cw[303] ^ cw[305] ^ cw[307] ^ cw[309] ^ cw[311] ^ cw[313] ^ cw[315] ^ cw[317] ^ cw[319] ^ cw[321] ^ cw[323] ^ cw[325] ^ cw[327] ^ cw[329] ^ cw[331] ^ cw[333] ^ cw[335] ^ cw[337] ^ cw[339] ^ cw[341] ^ cw[343] ^ cw[345] ^ cw[347] ^ cw[349] ^ cw[351] ^ cw[353] ^ cw[355] ^ cw[357] ^ cw[359] ^ cw[361] ^ cw[363] ^ cw[365] ^ cw[367] ^ cw[369] ^ cw[371] ^ cw[373] ^ cw[375] ^ cw[377] ^ cw[379] ^ cw[381] ^ cw[383] ^ cw[385] ^ cw[387] ^ cw[389] ^ cw[391] ^ cw[393] ^ cw[395] ^ cw[397] ^ cw[399] ^ cw[401] ^ cw[403] ^ cw[405] ^ cw[407] ^ cw[409] ^ cw[411] ^ cw[413] ^ cw[415] ^ cw[417] ^ cw[419] ^ cw[421] ^ cw[423] ^ cw[425] ^ cw[427] ^ cw[429] ^ cw[431] ^ cw[433] ^ cw[435] ^ cw[437] ^ cw[439] ^ cw[440] ^ cw[442] ^ cw[444] ^ cw[446] ^ cw[448] ^ cw[450] ^ cw[452] ^ cw[454] ^ cw[456] ^ cw[458] ^ cw[460] ^ cw[462] ^ cw[464] ^ cw[466] ^ cw[468] ^ cw[470] ^ cw[472] ^ cw[474] ^ cw[476] ^ cw[478] ^ cw[480] ^ cw[482] ^ cw[484] ^ cw[486] ^ cw[488] ^ cw[490] ^ cw[492] ^ cw[494] ^ cw[496] ^ cw[498] ^ cw[500] ^ cw[502] ^ cw[504] ^ cw[506] ^ cw[508] ^ cw[510] ^ cw[513] ^ cw[515] ^ cw[517] ^ cw[519] ^ cw[521] ^ cw[523] ^ cw[525] ^ cw[527] ^ cw[529] ^ cw[531] ^ cw[533] ^ cw[535] ^ cw[537] ^ cw[539] ^ cw[541] ^ cw[543] ^ cw[545] ^ cw[547] ^ cw[549] ^ cw[551] ^ cw[553] ^ cw[555] ^ cw[557] ^ cw[559] ^ cw[561] ^ cw[563] ^ cw[565] ^ cw[567] ^ cw[569] ^ cw[571] ^ cw[573] ^ cw[575] ^ cw[577] ^ cw[579] ^ cw[581] ^ cw[583] ^ cw[585] ^ cw[587] ^ cw[589] ^ cw[591] ^ cw[593] ^ cw[595] ^ cw[597] ^ cw[599] ^ cw[601] ^ cw[603] ^ cw[605] ^ cw[607] ^ cw[609] ^ cw[611] ^ cw[613] ^ cw[615] ^ cw[617] ^ cw[619] ^ cw[621] ^ cw[623] ^ cw[625] ^ cw[627] ^ cw[629] ^ cw[631] ^ cw[633] ^ cw[635] ^ cw[637] ^ cw[639] ^ cw[641] ^ cw[643] ^ cw[645] ^ cw[647] ^ cw[649] ^ cw[651] ^ cw[653] ^ cw[655] ^ cw[657] ^ cw[659] ^ cw[661] ^ cw[663] ^ cw[665] ^ cw[667] ^ cw[669] ^ cw[671] ^ cw[673] ^ cw[675] ^ cw[677] ^ cw[679] ^ cw[680] ^ cw[682] ^ cw[684] ^ cw[686] ^ cw[688] ^ cw[690] ^ cw[692] ^ cw[694] ^ cw[696] ^ cw[698] ^ cw[700] ^ cw[702] ^ cw[704] ^ cw[706] ^ cw[708] ^ cw[710] ^ cw[712] ^ cw[714] ^ cw[716] ^ cw[718] ^ cw[720] ^ cw[722] ^ cw[724] ^ cw[726] ^ cw[728] ^ cw[730] ^ cw[732] ^ cw[734] ^ cw[736] ^ cw[738] ^ cw[740] ^ cw[742] ^ cw[744] ^ cw[746] ^ cw[748] ^ cw[750] ^ cw[752] ^ cw[754] ^ cw[756] ^ cw[758] ^ cw[760] ^ cw[762] ^ cw[764] ^ cw[766] ^ cw[768] ^ cw[770] ^ cw[772] ^ cw[774] ^ cw[776] ^ cw[778] ^ cw[780] ^ cw[782] ^ cw[784] ^ cw[786] ^ cw[788] ^ cw[790] ^ cw[792] ^ cw[794] ^ cw[796] ^ cw[798] ^ cw[800] ^ cw[802] ^ cw[804] ^ cw[806] ^ cw[808] ^ cw[810] ^ cw[812] ^ cw[814] ^ cw[816] ^ cw[818] ^ cw[820] ^ cw[822] ^ cw[824] ^ cw[826] ^ cw[828] ^ cw[830] ^ cw[832] ^ cw[834] ^ cw[836] ^ cw[838] ^ cw[840] ^ cw[842] ^ cw[844] ^ cw[846] ^ cw[849] ^ cw[851] ^ cw[853] ^ cw[855] ^ cw[857] ^ cw[859] ^ cw[861] ^ cw[863] ^ cw[865] ^ cw[867] ^ cw[869] ^ cw[871] ^ cw[873] ^ cw[875] ^ cw[877] ^ cw[879] ^ cw[881] ^ cw[883] ^ cw[885] ^ cw[887] ^ cw[889] ^ cw[891] ^ cw[893] ^ cw[895] ^ cw[897] ^ cw[899] ^ cw[901] ^ cw[903] ^ cw[905] ^ cw[907] ^ cw[909] ^ cw[911] ^ cw[913] ^ cw[915] ^ cw[917] ^ cw[919] ^ cw[921] ^ cw[923] ^ cw[925] ^ cw[927] ^ cw[929] ^ cw[931] ^ cw[933] ^ cw[935] ^ cw[937] ^ cw[939] ^ cw[941] ^ cw[943] ^ cw[945] ^ cw[947] ^ cw[949] ^ cw[951] ^ cw[953] ^ cw[955] ^ cw[957] ^ cw[959] ^ cw[961] ^ cw[963] ^ cw[965] ^ cw[967] ^ cw[969] ^ cw[971] ^ cw[973] ^ cw[975] ^ cw[977] ^ cw[979] ^ cw[981] ^ cw[983] ^ cw[985] ^ cw[987] ^ cw[989] ^ cw[991] ^ cw[993] ^ cw[995] ^ cw[997] ^ cw[999] ^ cw[1001] ^ cw[1003] ^ cw[1005] ^ cw[1007] ^ cw[1009] ^ cw[1011] ^ cw[1013] ^ cw[1015] ^ cw[1017] ^ cw[1019] ^ cw[1021] ^ cw[1023] ^ cw[1025] ^ cw[1027] ^ cw[1029] ^ cw[1031] ^ cw[1033] ^ cw[1035] ^ cw[1037] ^ cw[1039] ^ cw[1041] ^ cw[1043] ^ cw[1045] ^ cw[1047] ^ cw[1049] ^ cw[1051] ^ cw[1053] ^ cw[1055] ^ cw[1057] ^ cw[1059] ^ cw[1061] ^ cw[1063] ^ cw[1065] ^ cw[1067] ^ cw[1069] ^ cw[1071] ^ cw[1073] ^ cw[1075] ^ cw[1077] ^ cw[1079] ^ cw[1081] ^ cw[1083] ^ cw[1085] ^ cw[1087] ^ cw[1089] ^ cw[1091] ^ cw[1093] ^ cw[1095] ^ cw[1097] ^ cw[1099] ^ cw[1100] ^ cw[1102] ^ cw[1104] ^ cw[1106] ^ cw[1108] ^ cw[1110] ^ cw[1112] ^ cw[1114] ^ cw[1116] ^ cw[1118] ^ cw[1120] ^ cw[1122] ^ cw[1124] ^ cw[1126] ^ cw[1128] ^ cw[1130] ^ cw[1132] ^ cw[1134] ^ cw[1136] ^ cw[1138] ^ cw[1140] ^ cw[1142] ^ cw[1144] ^ cw[1146] ^ cw[1148] ^ cw[1150] ^ cw[1152] ^ cw[1154] ^ cw[1156] ^ cw[1158] ^ cw[1160] ^ cw[1162] ^ cw[1164] ^ cw[1166] ^ cw[1168] ^ cw[1170] ^ cw[1172] ^ cw[1174] ^ cw[1176] ^ cw[1178] ^ cw[1180] ^ cw[1182] ^ cw[1184] ^ cw[1186] ^ cw[1188] ^ cw[1190] ^ cw[1192] ^ cw[1194] ^ cw[1196] ^ cw[1198] ^ cw[1200] ^ cw[1202] ^ cw[1204] ^ cw[1206] ^ cw[1208] ^ cw[1210] ^ cw[1212] ^ cw[1214] ^ cw[1216] ^ cw[1218] ^ cw[1220] ^ cw[1222] ^ cw[1224] ^ cw[1226] ^ cw[1228] ^ cw[1230] ^ cw[1232] ^ cw[1234] ^ cw[1236] ^ cw[1238] ^ cw[1240] ^ cw[1242] ^ cw[1244] ^ cw[1246] ^ cw[1248] ^ cw[1250] ^ cw[1252] ^ cw[1254] ^ cw[1256] ^ cw[1258] ^ cw[1260] ^ cw[1262] ^ cw[1264] ^ cw[1266] ^ cw[1269] ^ cw[1271] ^ cw[1273] ^ cw[1275] ^ cw[1277] ^ cw[1279] ^ cw[1281] ^ cw[1283] ^ cw[1285] ^ cw[1287] ^ cw[1289] ^ cw[1291] ^ cw[1293] ^ cw[1295] ^ cw[1297] ^ cw[1299] ^ cw[1301] ^ cw[1303] ^ cw[1305] ^ cw[1307] ^ cw[1309] ^ cw[1311] ^ cw[1313] ^ cw[1315] ^ cw[1317] ^ cw[1319] ^ cw[1321] ^ cw[1323] ^ cw[1325] ^ cw[1327] ^ cw[1329] ^ cw[1331] ^ cw[1333] ^ cw[1335] ^ cw[1337] ^ cw[1339] ^ cw[1341] ^ cw[1343] ^ cw[1345] ^ cw[1347] ^ cw[1349] ^ cw[1351] ^ cw[1353] ^ cw[1355] ^ cw[1357] ^ cw[1359] ^ cw[1361] ^ cw[1363] ^ cw[1365] ^ cw[1367] ^ cw[1369] ^ cw[1371] ^ cw[1373] ^ cw[1375] ^ cw[1377] ^ cw[1379] ^ cw[1381] ^ cw[1383] ^ cw[1385] ^ cw[1387] ^ cw[1389] ^ cw[1391] ^ cw[1393] ^ cw[1395] ^ cw[1397] ^ cw[1399] ^ cw[1401] ^ cw[1403] ^ cw[1405] ^ cw[1407] ^ cw[1409] ^ cw[1411] ^ cw[1413] ^ cw[1415] ^ cw[1417] ^ cw[1419] ^ cw[1421] ^ cw[1423] ^ cw[1425] ^ cw[1427] ^ cw[1429] ^ cw[1431] ^ cw[1433] ^ cw[1435] ^ cw[1437] ^ cw[1439] ^ cw[1441] ^ cw[1443] ^ cw[1445] ^ cw[1447] ^ cw[1449] ^ cw[1451] ^ cw[1453] ^ cw[1455] ^ cw[1457] ^ cw[1459] ^ cw[1461] ^ cw[1463] ^ cw[1465] ^ cw[1467] ^ cw[1469] ^ cw[1471] ^ cw[1473] ^ cw[1475] ^ cw[1477] ^ cw[1479] ^ cw[1481] ^ cw[1483] ^ cw[1485] ^ cw[1487] ^ cw[1489] ^ cw[1491] ^ cw[1493] ^ cw[1495] ^ cw[1497] ^ cw[1499] ^ cw[1501] ^ cw[1503] ^ cw[1505] ^ cw[1507] ^ cw[1509] ^ cw[1511] ^ cw[1513] ^ cw[1515] ^ cw[1517] ^ cw[1519] ^ cw[1520] ^ cw[1522] ^ cw[1524] ^ cw[1526] ^ cw[1528] ^ cw[1530] ^ cw[1532] ^ cw[1534] ^ cw[1536] ^ cw[1538] ^ cw[1540] ^ cw[1542] ^ cw[1544] ^ cw[1546] ^ cw[1548] ^ cw[1550] ^ cw[1552] ^ cw[1554] ^ cw[1556] ^ cw[1558] ^ cw[1560] ^ cw[1562] ^ cw[1564] ^ cw[1566] ^ cw[1568] ^ cw[1570] ^ cw[1572] ^ cw[1574] ^ cw[1576] ^ cw[1578] ^ cw[1580] ^ cw[1582] ^ cw[1584] ^ cw[1586] ^ cw[1588] ^ cw[1590] ^ cw[1592] ^ cw[1594] ^ cw[1596] ^ cw[1598] ^ cw[1600] ^ cw[1602] ^ cw[1604] ^ cw[1606] ^ cw[1608] ^ cw[1610] ^ cw[1612] ^ cw[1614] ^ cw[1616] ^ cw[1618] ^ cw[1620] ^ cw[1622] ^ cw[1624] ^ cw[1626] ^ cw[1628] ^ cw[1630] ^ cw[1632] ^ cw[1634] ^ cw[1636] ^ cw[1638] ^ cw[1640] ^ cw[1642] ^ cw[1644] ^ cw[1646] ^ cw[1648] ^ cw[1650] ^ cw[1652] ^ cw[1654] ^ cw[1656] ^ cw[1658] ^ cw[1660] ^ cw[1662] ^ cw[1664] ^ cw[1666] ^ cw[1668] ^ cw[1670] ^ cw[1672] ^ cw[1674] ^ cw[1676] ^ cw[1678] ^ cw[1680] ^ cw[1682] ^ cw[1684] ^ cw[1686] ^ cw[1688] ^ cw[1690] ^ cw[1692] ^ cw[1694] ^ cw[1696] ^ cw[1698] ^ cw[1700] ^ cw[1702] ^ cw[1704] ^ cw[1706] ^ cw[1708] ^ cw[1710] ^ cw[1712] ^ cw[1714] ^ cw[1716] ^ cw[1718] ^ cw[1720] ^ cw[1722] ^ cw[1724] ^ cw[1726] ^ cw[1728] ^ cw[1730] ^ cw[1732] ^ cw[1734] ^ cw[1736] ^ cw[1738] ^ cw[1740] ^ cw[1742] ^ cw[1744] ^ cw[1746] ^ cw[1748] ^ cw[1750] ^ cw[1752] ^ cw[1754] ^ cw[1756] ^ cw[1758] ^ cw[1760] ^ cw[1762] ^ cw[1764] ^ cw[1766] ^ cw[1768] ^ cw[1770] ^ cw[1773] ^ cw[1775] ^ cw[1777] ^ cw[1779] ^ cw[1781] ^ cw[1783] ^ cw[1785] ^ cw[1787] ^ cw[1789] ^ cw[1791] ^ cw[1793] ^ cw[1795] ^ cw[1797] ^ cw[1799] ^ cw[1801] ^ cw[1803] ^ cw[1805] ^ cw[1807] ^ cw[1809] ^ cw[1811] ^ cw[1813] ^ cw[1815] ^ cw[1817] ^ cw[1819] ^ cw[1821] ^ cw[1823] ^ cw[1825] ^ cw[1827] ^ cw[1829] ^ cw[1831] ^ cw[1833] ^ cw[1835] ^ cw[1837] ^ cw[1839] ^ cw[1841] ^ cw[1843] ^ cw[1845] ^ cw[1847] ^ cw[1849] ^ cw[1851] ^ cw[1853] ^ cw[1855] ^ cw[1857] ^ cw[1859] ^ cw[1861] ^ cw[1863] ^ cw[1865] ^ cw[1867] ^ cw[1869] ^ cw[1871] ^ cw[1873] ^ cw[1875] ^ cw[1877] ^ cw[1879] ^ cw[1881] ^ cw[1883] ^ cw[1885] ^ cw[1887] ^ cw[1889] ^ cw[1891] ^ cw[1893] ^ cw[1895] ^ cw[1897] ^ cw[1899] ^ cw[1901] ^ cw[1903] ^ cw[1905] ^ cw[1907] ^ cw[1909] ^ cw[1911] ^ cw[1913] ^ cw[1915] ^ cw[1917] ^ cw[1919] ^ cw[1921] ^ cw[1923] ^ cw[1925] ^ cw[1927] ^ cw[1929] ^ cw[1931] ^ cw[1933] ^ cw[1935] ^ cw[1937] ^ cw[1939] ^ cw[1941] ^ cw[1943] ^ cw[1945] ^ cw[1947] ^ cw[1949] ^ cw[1951] ^ cw[1953] ^ cw[1955] ^ cw[1957] ^ cw[1959] ^ cw[1961] ^ cw[1963] ^ cw[1965] ^ cw[1967] ^ cw[1969] ^ cw[1971] ^ cw[1973] ^ cw[1975] ^ cw[1977] ^ cw[1979] ^ cw[1981] ^ cw[1983] ^ cw[1985] ^ cw[1987] ^ cw[1989] ^ cw[1991] ^ cw[1993] ^ cw[1995] ^ cw[1997] ^ cw[1999] ^ cw[2001] ^ cw[2003] ^ cw[2005] ^ cw[2007] ^ cw[2009] ^ cw[2011] ^ cw[2013] ^ cw[2015] ^ cw[2017] ^ cw[2019] ^ cw[2021] ^ cw[2023] ^ cw[2024] ^ cw[2025] ^ cw[2026] ^ cw[2027] ^ cw[2028] ^ cw[2029] ^ cw[2030] ^ cw[2031] ^ cw[2032] ^ cw[2034] ^ cw[2035] ^ cw[2045];
    assign syndrome[1] = cw[0] ^ cw[2] ^ cw[4] ^ cw[6] ^ cw[8] ^ cw[10] ^ cw[12] ^ cw[14] ^ cw[16] ^ cw[18] ^ cw[21] ^ cw[23] ^ cw[25] ^ cw[27] ^ cw[29] ^ cw[31] ^ cw[33] ^ cw[35] ^ cw[37] ^ cw[39] ^ cw[41] ^ cw[43] ^ cw[45] ^ cw[47] ^ cw[49] ^ cw[51] ^ cw[53] ^ cw[55] ^ cw[57] ^ cw[59] ^ cw[61] ^ cw[63] ^ cw[65] ^ cw[67] ^ cw[69] ^ cw[71] ^ cw[73] ^ cw[75] ^ cw[77] ^ cw[79] ^ cw[81] ^ cw[83] ^ cw[85] ^ cw[87] ^ cw[89] ^ cw[91] ^ cw[93] ^ cw[95] ^ cw[97] ^ cw[99] ^ cw[101] ^ cw[103] ^ cw[105] ^ cw[107] ^ cw[109] ^ cw[110] ^ cw[112] ^ cw[114] ^ cw[116] ^ cw[118] ^ cw[120] ^ cw[122] ^ cw[124] ^ cw[126] ^ cw[128] ^ cw[130] ^ cw[132] ^ cw[134] ^ cw[136] ^ cw[138] ^ cw[140] ^ cw[142] ^ cw[144] ^ cw[146] ^ cw[148] ^ cw[150] ^ cw[152] ^ cw[154] ^ cw[156] ^ cw[158] ^ cw[160] ^ cw[162] ^ cw[164] ^ cw[166] ^ cw[168] ^ cw[170] ^ cw[172] ^ cw[174] ^ cw[176] ^ cw[178] ^ cw[180] ^ cw[182] ^ cw[184] ^ cw[186] ^ cw[188] ^ cw[190] ^ cw[192] ^ cw[194] ^ cw[196] ^ cw[198] ^ cw[201] ^ cw[203] ^ cw[205] ^ cw[207] ^ cw[209] ^ cw[211] ^ cw[213] ^ cw[215] ^ cw[217] ^ cw[219] ^ cw[221] ^ cw[223] ^ cw[225] ^ cw[227] ^ cw[229] ^ cw[231] ^ cw[233] ^ cw[235] ^ cw[237] ^ cw[239] ^ cw[241] ^ cw[243] ^ cw[245] ^ cw[247] ^ cw[249] ^ cw[251] ^ cw[253] ^ cw[255] ^ cw[257] ^ cw[259] ^ cw[261] ^ cw[263] ^ cw[265] ^ cw[267] ^ cw[269] ^ cw[271] ^ cw[273] ^ cw[275] ^ cw[277] ^ cw[279] ^ cw[281] ^ cw[283] ^ cw[285] ^ cw[287] ^ cw[289] ^ cw[291] ^ cw[293] ^ cw[295] ^ cw[297] ^ cw[299] ^ cw[301] ^ cw[303] ^ cw[305] ^ cw[307] ^ cw[309] ^ cw[311] ^ cw[313] ^ cw[315] ^ cw[317] ^ cw[319] ^ cw[321] ^ cw[323] ^ cw[325] ^ cw[327] ^ cw[329] ^ cw[331] ^ cw[333] ^ cw[335] ^ cw[337] ^ cw[339] ^ cw[341] ^ cw[343] ^ cw[345] ^ cw[347] ^ cw[349] ^ cw[351] ^ cw[353] ^ cw[355] ^ cw[357] ^ cw[359] ^ cw[361] ^ cw[363] ^ cw[365] ^ cw[367] ^ cw[369] ^ cw[371] ^ cw[373] ^ cw[375] ^ cw[377] ^ cw[379] ^ cw[381] ^ cw[383] ^ cw[385] ^ cw[387] ^ cw[389] ^ cw[391] ^ cw[393] ^ cw[395] ^ cw[397] ^ cw[399] ^ cw[401] ^ cw[403] ^ cw[405] ^ cw[407] ^ cw[409] ^ cw[411] ^ cw[413] ^ cw[415] ^ cw[417] ^ cw[419] ^ cw[421] ^ cw[423] ^ cw[425] ^ cw[427] ^ cw[429] ^ cw[431] ^ cw[433] ^ cw[435] ^ cw[437] ^ cw[439] ^ cw[440] ^ cw[442] ^ cw[444] ^ cw[446] ^ cw[448] ^ cw[450] ^ cw[452] ^ cw[454] ^ cw[456] ^ cw[458] ^ cw[460] ^ cw[462] ^ cw[464] ^ cw[466] ^ cw[468] ^ cw[470] ^ cw[472] ^ cw[474] ^ cw[476] ^ cw[478] ^ cw[480] ^ cw[482] ^ cw[484] ^ cw[486] ^ cw[488] ^ cw[490] ^ cw[492] ^ cw[494] ^ cw[496] ^ cw[498] ^ cw[500] ^ cw[502] ^ cw[504] ^ cw[506] ^ cw[508] ^ cw[510] ^ cw[512] ^ cw[514] ^ cw[516] ^ cw[518] ^ cw[520] ^ cw[522] ^ cw[524] ^ cw[526] ^ cw[528] ^ cw[530] ^ cw[532] ^ cw[534] ^ cw[536] ^ cw[538] ^ cw[540] ^ cw[542] ^ cw[544] ^ cw[546] ^ cw[548] ^ cw[550] ^ cw[552] ^ cw[554] ^ cw[556] ^ cw[558] ^ cw[560] ^ cw[562] ^ cw[564] ^ cw[566] ^ cw[568] ^ cw[570] ^ cw[572] ^ cw[574] ^ cw[576] ^ cw[578] ^ cw[580] ^ cw[582] ^ cw[584] ^ cw[586] ^ cw[588] ^ cw[590] ^ cw[592] ^ cw[594] ^ cw[596] ^ cw[598] ^ cw[600] ^ cw[602] ^ cw[604] ^ cw[606] ^ cw[608] ^ cw[610] ^ cw[612] ^ cw[614] ^ cw[616] ^ cw[618] ^ cw[620] ^ cw[622] ^ cw[624] ^ cw[626] ^ cw[628] ^ cw[630] ^ cw[632] ^ cw[634] ^ cw[636] ^ cw[638] ^ cw[640] ^ cw[642] ^ cw[644] ^ cw[646] ^ cw[648] ^ cw[650] ^ cw[652] ^ cw[654] ^ cw[656] ^ cw[658] ^ cw[660] ^ cw[662] ^ cw[664] ^ cw[666] ^ cw[668] ^ cw[670] ^ cw[672] ^ cw[674] ^ cw[676] ^ cw[678] ^ cw[681] ^ cw[683] ^ cw[685] ^ cw[687] ^ cw[689] ^ cw[691] ^ cw[693] ^ cw[695] ^ cw[697] ^ cw[699] ^ cw[701] ^ cw[703] ^ cw[705] ^ cw[707] ^ cw[709] ^ cw[711] ^ cw[713] ^ cw[715] ^ cw[717] ^ cw[719] ^ cw[721] ^ cw[723] ^ cw[725] ^ cw[727] ^ cw[729] ^ cw[731] ^ cw[733] ^ cw[735] ^ cw[737] ^ cw[739] ^ cw[741] ^ cw[743] ^ cw[745] ^ cw[747] ^ cw[749] ^ cw[751] ^ cw[753] ^ cw[755] ^ cw[757] ^ cw[759] ^ cw[761] ^ cw[763] ^ cw[765] ^ cw[767] ^ cw[769] ^ cw[771] ^ cw[773] ^ cw[775] ^ cw[777] ^ cw[779] ^ cw[781] ^ cw[783] ^ cw[785] ^ cw[787] ^ cw[789] ^ cw[791] ^ cw[793] ^ cw[795] ^ cw[797] ^ cw[799] ^ cw[801] ^ cw[803] ^ cw[805] ^ cw[807] ^ cw[809] ^ cw[811] ^ cw[813] ^ cw[815] ^ cw[817] ^ cw[819] ^ cw[821] ^ cw[823] ^ cw[825] ^ cw[827] ^ cw[829] ^ cw[831] ^ cw[833] ^ cw[835] ^ cw[837] ^ cw[839] ^ cw[841] ^ cw[843] ^ cw[845] ^ cw[847] ^ cw[849] ^ cw[851] ^ cw[853] ^ cw[855] ^ cw[857] ^ cw[859] ^ cw[861] ^ cw[863] ^ cw[865] ^ cw[867] ^ cw[869] ^ cw[871] ^ cw[873] ^ cw[875] ^ cw[877] ^ cw[879] ^ cw[881] ^ cw[883] ^ cw[885] ^ cw[887] ^ cw[889] ^ cw[891] ^ cw[893] ^ cw[895] ^ cw[897] ^ cw[899] ^ cw[901] ^ cw[903] ^ cw[905] ^ cw[907] ^ cw[909] ^ cw[911] ^ cw[913] ^ cw[915] ^ cw[917] ^ cw[919] ^ cw[921] ^ cw[923] ^ cw[925] ^ cw[927] ^ cw[929] ^ cw[931] ^ cw[933] ^ cw[935] ^ cw[937] ^ cw[939] ^ cw[941] ^ cw[943] ^ cw[945] ^ cw[947] ^ cw[949] ^ cw[951] ^ cw[953] ^ cw[955] ^ cw[957] ^ cw[959] ^ cw[961] ^ cw[963] ^ cw[965] ^ cw[967] ^ cw[969] ^ cw[971] ^ cw[973] ^ cw[975] ^ cw[977] ^ cw[979] ^ cw[981] ^ cw[983] ^ cw[985] ^ cw[987] ^ cw[989] ^ cw[991] ^ cw[993] ^ cw[995] ^ cw[997] ^ cw[999] ^ cw[1001] ^ cw[1003] ^ cw[1005] ^ cw[1007] ^ cw[1009] ^ cw[1011] ^ cw[1013] ^ cw[1015] ^ cw[1017] ^ cw[1019] ^ cw[1021] ^ cw[1023] ^ cw[1025] ^ cw[1027] ^ cw[1029] ^ cw[1031] ^ cw[1033] ^ cw[1035] ^ cw[1037] ^ cw[1039] ^ cw[1041] ^ cw[1043] ^ cw[1045] ^ cw[1047] ^ cw[1049] ^ cw[1051] ^ cw[1053] ^ cw[1055] ^ cw[1057] ^ cw[1059] ^ cw[1061] ^ cw[1063] ^ cw[1065] ^ cw[1067] ^ cw[1069] ^ cw[1071] ^ cw[1073] ^ cw[1075] ^ cw[1077] ^ cw[1079] ^ cw[1081] ^ cw[1083] ^ cw[1085] ^ cw[1087] ^ cw[1089] ^ cw[1091] ^ cw[1093] ^ cw[1095] ^ cw[1097] ^ cw[1099] ^ cw[1100] ^ cw[1102] ^ cw[1104] ^ cw[1106] ^ cw[1108] ^ cw[1110] ^ cw[1112] ^ cw[1114] ^ cw[1116] ^ cw[1118] ^ cw[1120] ^ cw[1122] ^ cw[1124] ^ cw[1126] ^ cw[1128] ^ cw[1130] ^ cw[1132] ^ cw[1134] ^ cw[1136] ^ cw[1138] ^ cw[1140] ^ cw[1142] ^ cw[1144] ^ cw[1146] ^ cw[1148] ^ cw[1150] ^ cw[1152] ^ cw[1154] ^ cw[1156] ^ cw[1158] ^ cw[1160] ^ cw[1162] ^ cw[1164] ^ cw[1166] ^ cw[1168] ^ cw[1170] ^ cw[1172] ^ cw[1174] ^ cw[1176] ^ cw[1178] ^ cw[1180] ^ cw[1182] ^ cw[1184] ^ cw[1186] ^ cw[1188] ^ cw[1190] ^ cw[1192] ^ cw[1194] ^ cw[1196] ^ cw[1198] ^ cw[1200] ^ cw[1202] ^ cw[1204] ^ cw[1206] ^ cw[1208] ^ cw[1210] ^ cw[1212] ^ cw[1214] ^ cw[1216] ^ cw[1218] ^ cw[1220] ^ cw[1222] ^ cw[1224] ^ cw[1226] ^ cw[1228] ^ cw[1230] ^ cw[1232] ^ cw[1234] ^ cw[1236] ^ cw[1238] ^ cw[1240] ^ cw[1242] ^ cw[1244] ^ cw[1246] ^ cw[1248] ^ cw[1250] ^ cw[1252] ^ cw[1254] ^ cw[1256] ^ cw[1258] ^ cw[1260] ^ cw[1262] ^ cw[1264] ^ cw[1266] ^ cw[1268] ^ cw[1270] ^ cw[1272] ^ cw[1274] ^ cw[1276] ^ cw[1278] ^ cw[1280] ^ cw[1282] ^ cw[1284] ^ cw[1286] ^ cw[1288] ^ cw[1290] ^ cw[1292] ^ cw[1294] ^ cw[1296] ^ cw[1298] ^ cw[1300] ^ cw[1302] ^ cw[1304] ^ cw[1306] ^ cw[1308] ^ cw[1310] ^ cw[1312] ^ cw[1314] ^ cw[1316] ^ cw[1318] ^ cw[1320] ^ cw[1322] ^ cw[1324] ^ cw[1326] ^ cw[1328] ^ cw[1330] ^ cw[1332] ^ cw[1334] ^ cw[1336] ^ cw[1338] ^ cw[1340] ^ cw[1342] ^ cw[1344] ^ cw[1346] ^ cw[1348] ^ cw[1350] ^ cw[1352] ^ cw[1354] ^ cw[1356] ^ cw[1358] ^ cw[1360] ^ cw[1362] ^ cw[1364] ^ cw[1366] ^ cw[1368] ^ cw[1370] ^ cw[1372] ^ cw[1374] ^ cw[1376] ^ cw[1378] ^ cw[1380] ^ cw[1382] ^ cw[1384] ^ cw[1386] ^ cw[1388] ^ cw[1390] ^ cw[1392] ^ cw[1394] ^ cw[1396] ^ cw[1398] ^ cw[1400] ^ cw[1402] ^ cw[1404] ^ cw[1406] ^ cw[1408] ^ cw[1410] ^ cw[1412] ^ cw[1414] ^ cw[1416] ^ cw[1418] ^ cw[1420] ^ cw[1422] ^ cw[1424] ^ cw[1426] ^ cw[1428] ^ cw[1430] ^ cw[1432] ^ cw[1434] ^ cw[1436] ^ cw[1438] ^ cw[1440] ^ cw[1442] ^ cw[1444] ^ cw[1446] ^ cw[1448] ^ cw[1450] ^ cw[1452] ^ cw[1454] ^ cw[1456] ^ cw[1458] ^ cw[1460] ^ cw[1462] ^ cw[1464] ^ cw[1466] ^ cw[1468] ^ cw[1470] ^ cw[1472] ^ cw[1474] ^ cw[1476] ^ cw[1478] ^ cw[1480] ^ cw[1482] ^ cw[1484] ^ cw[1486] ^ cw[1488] ^ cw[1490] ^ cw[1492] ^ cw[1494] ^ cw[1496] ^ cw[1498] ^ cw[1500] ^ cw[1502] ^ cw[1504] ^ cw[1506] ^ cw[1508] ^ cw[1510] ^ cw[1512] ^ cw[1514] ^ cw[1516] ^ cw[1518] ^ cw[1521] ^ cw[1523] ^ cw[1525] ^ cw[1527] ^ cw[1529] ^ cw[1531] ^ cw[1533] ^ cw[1535] ^ cw[1537] ^ cw[1539] ^ cw[1541] ^ cw[1543] ^ cw[1545] ^ cw[1547] ^ cw[1549] ^ cw[1551] ^ cw[1553] ^ cw[1555] ^ cw[1557] ^ cw[1559] ^ cw[1561] ^ cw[1563] ^ cw[1565] ^ cw[1567] ^ cw[1569] ^ cw[1571] ^ cw[1573] ^ cw[1575] ^ cw[1577] ^ cw[1579] ^ cw[1581] ^ cw[1583] ^ cw[1585] ^ cw[1587] ^ cw[1589] ^ cw[1591] ^ cw[1593] ^ cw[1595] ^ cw[1597] ^ cw[1599] ^ cw[1601] ^ cw[1603] ^ cw[1605] ^ cw[1607] ^ cw[1609] ^ cw[1611] ^ cw[1613] ^ cw[1615] ^ cw[1617] ^ cw[1619] ^ cw[1621] ^ cw[1623] ^ cw[1625] ^ cw[1627] ^ cw[1629] ^ cw[1631] ^ cw[1633] ^ cw[1635] ^ cw[1637] ^ cw[1639] ^ cw[1641] ^ cw[1643] ^ cw[1645] ^ cw[1647] ^ cw[1649] ^ cw[1651] ^ cw[1653] ^ cw[1655] ^ cw[1657] ^ cw[1659] ^ cw[1661] ^ cw[1663] ^ cw[1665] ^ cw[1667] ^ cw[1669] ^ cw[1671] ^ cw[1673] ^ cw[1675] ^ cw[1677] ^ cw[1679] ^ cw[1681] ^ cw[1683] ^ cw[1685] ^ cw[1687] ^ cw[1689] ^ cw[1691] ^ cw[1693] ^ cw[1695] ^ cw[1697] ^ cw[1699] ^ cw[1701] ^ cw[1703] ^ cw[1705] ^ cw[1707] ^ cw[1709] ^ cw[1711] ^ cw[1713] ^ cw[1715] ^ cw[1717] ^ cw[1719] ^ cw[1721] ^ cw[1723] ^ cw[1725] ^ cw[1727] ^ cw[1729] ^ cw[1731] ^ cw[1733] ^ cw[1735] ^ cw[1737] ^ cw[1739] ^ cw[1741] ^ cw[1743] ^ cw[1745] ^ cw[1747] ^ cw[1749] ^ cw[1751] ^ cw[1753] ^ cw[1755] ^ cw[1757] ^ cw[1759] ^ cw[1761] ^ cw[1763] ^ cw[1765] ^ cw[1767] ^ cw[1769] ^ cw[1771] ^ cw[1773] ^ cw[1775] ^ cw[1777] ^ cw[1779] ^ cw[1781] ^ cw[1783] ^ cw[1785] ^ cw[1787] ^ cw[1789] ^ cw[1791] ^ cw[1793] ^ cw[1795] ^ cw[1797] ^ cw[1799] ^ cw[1801] ^ cw[1803] ^ cw[1805] ^ cw[1807] ^ cw[1809] ^ cw[1811] ^ cw[1813] ^ cw[1815] ^ cw[1817] ^ cw[1819] ^ cw[1821] ^ cw[1823] ^ cw[1825] ^ cw[1827] ^ cw[1829] ^ cw[1831] ^ cw[1833] ^ cw[1835] ^ cw[1837] ^ cw[1839] ^ cw[1841] ^ cw[1843] ^ cw[1845] ^ cw[1847] ^ cw[1849] ^ cw[1851] ^ cw[1853] ^ cw[1855] ^ cw[1857] ^ cw[1859] ^ cw[1861] ^ cw[1863] ^ cw[1865] ^ cw[1867] ^ cw[1869] ^ cw[1871] ^ cw[1873] ^ cw[1875] ^ cw[1877] ^ cw[1879] ^ cw[1881] ^ cw[1883] ^ cw[1885] ^ cw[1887] ^ cw[1889] ^ cw[1891] ^ cw[1893] ^ cw[1895] ^ cw[1897] ^ cw[1899] ^ cw[1901] ^ cw[1903] ^ cw[1905] ^ cw[1907] ^ cw[1909] ^ cw[1911] ^ cw[1913] ^ cw[1915] ^ cw[1917] ^ cw[1919] ^ cw[1921] ^ cw[1923] ^ cw[1925] ^ cw[1927] ^ cw[1929] ^ cw[1931] ^ cw[1933] ^ cw[1935] ^ cw[1937] ^ cw[1939] ^ cw[1941] ^ cw[1943] ^ cw[1945] ^ cw[1947] ^ cw[1949] ^ cw[1951] ^ cw[1953] ^ cw[1955] ^ cw[1957] ^ cw[1959] ^ cw[1961] ^ cw[1963] ^ cw[1965] ^ cw[1967] ^ cw[1969] ^ cw[1971] ^ cw[1973] ^ cw[1975] ^ cw[1977] ^ cw[1979] ^ cw[1981] ^ cw[1983] ^ cw[1985] ^ cw[1987] ^ cw[1989] ^ cw[1991] ^ cw[1993] ^ cw[1995] ^ cw[1997] ^ cw[1999] ^ cw[2001] ^ cw[2003] ^ cw[2005] ^ cw[2007] ^ cw[2009] ^ cw[2011] ^ cw[2013] ^ cw[2015] ^ cw[2017] ^ cw[2019] ^ cw[2021] ^ cw[2023] ^ cw[2024] ^ cw[2025] ^ cw[2026] ^ cw[2027] ^ cw[2028] ^ cw[2029] ^ cw[2030] ^ cw[2031] ^ cw[2032] ^ cw[2033] ^ cw[2035] ^ cw[2046];
    assign syndrome[0] = cw[0] ^ cw[2] ^ cw[4] ^ cw[6] ^ cw[8] ^ cw[10] ^ cw[12] ^ cw[14] ^ cw[16] ^ cw[18] ^ cw[20] ^ cw[22] ^ cw[24] ^ cw[26] ^ cw[28] ^ cw[30] ^ cw[32] ^ cw[34] ^ cw[36] ^ cw[38] ^ cw[40] ^ cw[42] ^ cw[44] ^ cw[46] ^ cw[48] ^ cw[50] ^ cw[52] ^ cw[54] ^ cw[56] ^ cw[58] ^ cw[60] ^ cw[62] ^ cw[64] ^ cw[66] ^ cw[68] ^ cw[70] ^ cw[72] ^ cw[74] ^ cw[76] ^ cw[78] ^ cw[80] ^ cw[82] ^ cw[84] ^ cw[86] ^ cw[88] ^ cw[90] ^ cw[92] ^ cw[94] ^ cw[96] ^ cw[98] ^ cw[100] ^ cw[102] ^ cw[104] ^ cw[106] ^ cw[108] ^ cw[111] ^ cw[113] ^ cw[115] ^ cw[117] ^ cw[119] ^ cw[121] ^ cw[123] ^ cw[125] ^ cw[127] ^ cw[129] ^ cw[131] ^ cw[133] ^ cw[135] ^ cw[137] ^ cw[139] ^ cw[141] ^ cw[143] ^ cw[145] ^ cw[147] ^ cw[149] ^ cw[151] ^ cw[153] ^ cw[155] ^ cw[157] ^ cw[159] ^ cw[161] ^ cw[163] ^ cw[165] ^ cw[167] ^ cw[169] ^ cw[171] ^ cw[173] ^ cw[175] ^ cw[177] ^ cw[179] ^ cw[181] ^ cw[183] ^ cw[185] ^ cw[187] ^ cw[189] ^ cw[191] ^ cw[193] ^ cw[195] ^ cw[197] ^ cw[199] ^ cw[201] ^ cw[203] ^ cw[205] ^ cw[207] ^ cw[209] ^ cw[211] ^ cw[213] ^ cw[215] ^ cw[217] ^ cw[219] ^ cw[221] ^ cw[223] ^ cw[225] ^ cw[227] ^ cw[229] ^ cw[231] ^ cw[233] ^ cw[235] ^ cw[237] ^ cw[239] ^ cw[241] ^ cw[243] ^ cw[245] ^ cw[247] ^ cw[249] ^ cw[251] ^ cw[253] ^ cw[255] ^ cw[257] ^ cw[259] ^ cw[261] ^ cw[263] ^ cw[265] ^ cw[267] ^ cw[269] ^ cw[271] ^ cw[273] ^ cw[275] ^ cw[277] ^ cw[279] ^ cw[281] ^ cw[283] ^ cw[285] ^ cw[287] ^ cw[289] ^ cw[291] ^ cw[293] ^ cw[295] ^ cw[297] ^ cw[299] ^ cw[301] ^ cw[303] ^ cw[305] ^ cw[307] ^ cw[309] ^ cw[311] ^ cw[313] ^ cw[315] ^ cw[317] ^ cw[319] ^ cw[321] ^ cw[323] ^ cw[325] ^ cw[327] ^ cw[329] ^ cw[331] ^ cw[333] ^ cw[335] ^ cw[337] ^ cw[339] ^ cw[341] ^ cw[343] ^ cw[345] ^ cw[347] ^ cw[349] ^ cw[351] ^ cw[353] ^ cw[355] ^ cw[357] ^ cw[359] ^ cw[361] ^ cw[363] ^ cw[365] ^ cw[367] ^ cw[369] ^ cw[371] ^ cw[373] ^ cw[375] ^ cw[377] ^ cw[379] ^ cw[381] ^ cw[383] ^ cw[385] ^ cw[387] ^ cw[389] ^ cw[391] ^ cw[393] ^ cw[395] ^ cw[397] ^ cw[399] ^ cw[401] ^ cw[403] ^ cw[405] ^ cw[407] ^ cw[409] ^ cw[411] ^ cw[413] ^ cw[415] ^ cw[417] ^ cw[419] ^ cw[421] ^ cw[423] ^ cw[425] ^ cw[427] ^ cw[429] ^ cw[431] ^ cw[433] ^ cw[435] ^ cw[437] ^ cw[439] ^ cw[440] ^ cw[442] ^ cw[444] ^ cw[446] ^ cw[448] ^ cw[450] ^ cw[452] ^ cw[454] ^ cw[456] ^ cw[458] ^ cw[460] ^ cw[462] ^ cw[464] ^ cw[466] ^ cw[468] ^ cw[470] ^ cw[472] ^ cw[474] ^ cw[476] ^ cw[478] ^ cw[480] ^ cw[482] ^ cw[484] ^ cw[486] ^ cw[488] ^ cw[490] ^ cw[492] ^ cw[494] ^ cw[496] ^ cw[498] ^ cw[500] ^ cw[502] ^ cw[504] ^ cw[506] ^ cw[508] ^ cw[510] ^ cw[512] ^ cw[514] ^ cw[516] ^ cw[518] ^ cw[520] ^ cw[522] ^ cw[524] ^ cw[526] ^ cw[528] ^ cw[530] ^ cw[532] ^ cw[534] ^ cw[536] ^ cw[538] ^ cw[540] ^ cw[542] ^ cw[544] ^ cw[546] ^ cw[548] ^ cw[550] ^ cw[552] ^ cw[554] ^ cw[556] ^ cw[558] ^ cw[560] ^ cw[562] ^ cw[564] ^ cw[566] ^ cw[568] ^ cw[570] ^ cw[572] ^ cw[574] ^ cw[576] ^ cw[578] ^ cw[580] ^ cw[582] ^ cw[584] ^ cw[586] ^ cw[588] ^ cw[590] ^ cw[592] ^ cw[594] ^ cw[596] ^ cw[598] ^ cw[600] ^ cw[602] ^ cw[604] ^ cw[606] ^ cw[608] ^ cw[610] ^ cw[612] ^ cw[614] ^ cw[616] ^ cw[618] ^ cw[620] ^ cw[622] ^ cw[624] ^ cw[626] ^ cw[628] ^ cw[630] ^ cw[632] ^ cw[634] ^ cw[636] ^ cw[638] ^ cw[640] ^ cw[642] ^ cw[644] ^ cw[646] ^ cw[648] ^ cw[650] ^ cw[652] ^ cw[654] ^ cw[656] ^ cw[658] ^ cw[660] ^ cw[662] ^ cw[664] ^ cw[666] ^ cw[668] ^ cw[670] ^ cw[672] ^ cw[674] ^ cw[676] ^ cw[678] ^ cw[680] ^ cw[682] ^ cw[684] ^ cw[686] ^ cw[688] ^ cw[690] ^ cw[692] ^ cw[694] ^ cw[696] ^ cw[698] ^ cw[700] ^ cw[702] ^ cw[704] ^ cw[706] ^ cw[708] ^ cw[710] ^ cw[712] ^ cw[714] ^ cw[716] ^ cw[718] ^ cw[720] ^ cw[722] ^ cw[724] ^ cw[726] ^ cw[728] ^ cw[730] ^ cw[732] ^ cw[734] ^ cw[736] ^ cw[738] ^ cw[740] ^ cw[742] ^ cw[744] ^ cw[746] ^ cw[748] ^ cw[750] ^ cw[752] ^ cw[754] ^ cw[756] ^ cw[758] ^ cw[760] ^ cw[762] ^ cw[764] ^ cw[766] ^ cw[768] ^ cw[770] ^ cw[772] ^ cw[774] ^ cw[776] ^ cw[778] ^ cw[780] ^ cw[782] ^ cw[784] ^ cw[786] ^ cw[788] ^ cw[790] ^ cw[792] ^ cw[794] ^ cw[796] ^ cw[798] ^ cw[800] ^ cw[802] ^ cw[804] ^ cw[806] ^ cw[808] ^ cw[810] ^ cw[812] ^ cw[814] ^ cw[816] ^ cw[818] ^ cw[820] ^ cw[822] ^ cw[824] ^ cw[826] ^ cw[828] ^ cw[830] ^ cw[832] ^ cw[834] ^ cw[836] ^ cw[838] ^ cw[840] ^ cw[842] ^ cw[844] ^ cw[846] ^ cw[848] ^ cw[850] ^ cw[852] ^ cw[854] ^ cw[856] ^ cw[858] ^ cw[860] ^ cw[862] ^ cw[864] ^ cw[866] ^ cw[868] ^ cw[870] ^ cw[872] ^ cw[874] ^ cw[876] ^ cw[878] ^ cw[880] ^ cw[882] ^ cw[884] ^ cw[886] ^ cw[888] ^ cw[890] ^ cw[892] ^ cw[894] ^ cw[896] ^ cw[898] ^ cw[900] ^ cw[902] ^ cw[904] ^ cw[906] ^ cw[908] ^ cw[910] ^ cw[912] ^ cw[914] ^ cw[916] ^ cw[918] ^ cw[920] ^ cw[922] ^ cw[924] ^ cw[926] ^ cw[928] ^ cw[930] ^ cw[932] ^ cw[934] ^ cw[936] ^ cw[938] ^ cw[940] ^ cw[942] ^ cw[944] ^ cw[946] ^ cw[948] ^ cw[950] ^ cw[952] ^ cw[954] ^ cw[956] ^ cw[958] ^ cw[960] ^ cw[962] ^ cw[964] ^ cw[966] ^ cw[968] ^ cw[970] ^ cw[972] ^ cw[974] ^ cw[976] ^ cw[978] ^ cw[980] ^ cw[982] ^ cw[984] ^ cw[986] ^ cw[988] ^ cw[990] ^ cw[992] ^ cw[994] ^ cw[996] ^ cw[998] ^ cw[1000] ^ cw[1002] ^ cw[1004] ^ cw[1006] ^ cw[1008] ^ cw[1010] ^ cw[1012] ^ cw[1014] ^ cw[1016] ^ cw[1018] ^ cw[1020] ^ cw[1022] ^ cw[1024] ^ cw[1026] ^ cw[1028] ^ cw[1030] ^ cw[1032] ^ cw[1034] ^ cw[1036] ^ cw[1038] ^ cw[1040] ^ cw[1042] ^ cw[1044] ^ cw[1046] ^ cw[1048] ^ cw[1050] ^ cw[1052] ^ cw[1054] ^ cw[1056] ^ cw[1058] ^ cw[1060] ^ cw[1062] ^ cw[1064] ^ cw[1066] ^ cw[1068] ^ cw[1070] ^ cw[1072] ^ cw[1074] ^ cw[1076] ^ cw[1078] ^ cw[1080] ^ cw[1082] ^ cw[1084] ^ cw[1086] ^ cw[1088] ^ cw[1090] ^ cw[1092] ^ cw[1094] ^ cw[1096] ^ cw[1098] ^ cw[1101] ^ cw[1103] ^ cw[1105] ^ cw[1107] ^ cw[1109] ^ cw[1111] ^ cw[1113] ^ cw[1115] ^ cw[1117] ^ cw[1119] ^ cw[1121] ^ cw[1123] ^ cw[1125] ^ cw[1127] ^ cw[1129] ^ cw[1131] ^ cw[1133] ^ cw[1135] ^ cw[1137] ^ cw[1139] ^ cw[1141] ^ cw[1143] ^ cw[1145] ^ cw[1147] ^ cw[1149] ^ cw[1151] ^ cw[1153] ^ cw[1155] ^ cw[1157] ^ cw[1159] ^ cw[1161] ^ cw[1163] ^ cw[1165] ^ cw[1167] ^ cw[1169] ^ cw[1171] ^ cw[1173] ^ cw[1175] ^ cw[1177] ^ cw[1179] ^ cw[1181] ^ cw[1183] ^ cw[1185] ^ cw[1187] ^ cw[1189] ^ cw[1191] ^ cw[1193] ^ cw[1195] ^ cw[1197] ^ cw[1199] ^ cw[1201] ^ cw[1203] ^ cw[1205] ^ cw[1207] ^ cw[1209] ^ cw[1211] ^ cw[1213] ^ cw[1215] ^ cw[1217] ^ cw[1219] ^ cw[1221] ^ cw[1223] ^ cw[1225] ^ cw[1227] ^ cw[1229] ^ cw[1231] ^ cw[1233] ^ cw[1235] ^ cw[1237] ^ cw[1239] ^ cw[1241] ^ cw[1243] ^ cw[1245] ^ cw[1247] ^ cw[1249] ^ cw[1251] ^ cw[1253] ^ cw[1255] ^ cw[1257] ^ cw[1259] ^ cw[1261] ^ cw[1263] ^ cw[1265] ^ cw[1267] ^ cw[1269] ^ cw[1271] ^ cw[1273] ^ cw[1275] ^ cw[1277] ^ cw[1279] ^ cw[1281] ^ cw[1283] ^ cw[1285] ^ cw[1287] ^ cw[1289] ^ cw[1291] ^ cw[1293] ^ cw[1295] ^ cw[1297] ^ cw[1299] ^ cw[1301] ^ cw[1303] ^ cw[1305] ^ cw[1307] ^ cw[1309] ^ cw[1311] ^ cw[1313] ^ cw[1315] ^ cw[1317] ^ cw[1319] ^ cw[1321] ^ cw[1323] ^ cw[1325] ^ cw[1327] ^ cw[1329] ^ cw[1331] ^ cw[1333] ^ cw[1335] ^ cw[1337] ^ cw[1339] ^ cw[1341] ^ cw[1343] ^ cw[1345] ^ cw[1347] ^ cw[1349] ^ cw[1351] ^ cw[1353] ^ cw[1355] ^ cw[1357] ^ cw[1359] ^ cw[1361] ^ cw[1363] ^ cw[1365] ^ cw[1367] ^ cw[1369] ^ cw[1371] ^ cw[1373] ^ cw[1375] ^ cw[1377] ^ cw[1379] ^ cw[1381] ^ cw[1383] ^ cw[1385] ^ cw[1387] ^ cw[1389] ^ cw[1391] ^ cw[1393] ^ cw[1395] ^ cw[1397] ^ cw[1399] ^ cw[1401] ^ cw[1403] ^ cw[1405] ^ cw[1407] ^ cw[1409] ^ cw[1411] ^ cw[1413] ^ cw[1415] ^ cw[1417] ^ cw[1419] ^ cw[1421] ^ cw[1423] ^ cw[1425] ^ cw[1427] ^ cw[1429] ^ cw[1431] ^ cw[1433] ^ cw[1435] ^ cw[1437] ^ cw[1439] ^ cw[1441] ^ cw[1443] ^ cw[1445] ^ cw[1447] ^ cw[1449] ^ cw[1451] ^ cw[1453] ^ cw[1455] ^ cw[1457] ^ cw[1459] ^ cw[1461] ^ cw[1463] ^ cw[1465] ^ cw[1467] ^ cw[1469] ^ cw[1471] ^ cw[1473] ^ cw[1475] ^ cw[1477] ^ cw[1479] ^ cw[1481] ^ cw[1483] ^ cw[1485] ^ cw[1487] ^ cw[1489] ^ cw[1491] ^ cw[1493] ^ cw[1495] ^ cw[1497] ^ cw[1499] ^ cw[1501] ^ cw[1503] ^ cw[1505] ^ cw[1507] ^ cw[1509] ^ cw[1511] ^ cw[1513] ^ cw[1515] ^ cw[1517] ^ cw[1519] ^ cw[1521] ^ cw[1523] ^ cw[1525] ^ cw[1527] ^ cw[1529] ^ cw[1531] ^ cw[1533] ^ cw[1535] ^ cw[1537] ^ cw[1539] ^ cw[1541] ^ cw[1543] ^ cw[1545] ^ cw[1547] ^ cw[1549] ^ cw[1551] ^ cw[1553] ^ cw[1555] ^ cw[1557] ^ cw[1559] ^ cw[1561] ^ cw[1563] ^ cw[1565] ^ cw[1567] ^ cw[1569] ^ cw[1571] ^ cw[1573] ^ cw[1575] ^ cw[1577] ^ cw[1579] ^ cw[1581] ^ cw[1583] ^ cw[1585] ^ cw[1587] ^ cw[1589] ^ cw[1591] ^ cw[1593] ^ cw[1595] ^ cw[1597] ^ cw[1599] ^ cw[1601] ^ cw[1603] ^ cw[1605] ^ cw[1607] ^ cw[1609] ^ cw[1611] ^ cw[1613] ^ cw[1615] ^ cw[1617] ^ cw[1619] ^ cw[1621] ^ cw[1623] ^ cw[1625] ^ cw[1627] ^ cw[1629] ^ cw[1631] ^ cw[1633] ^ cw[1635] ^ cw[1637] ^ cw[1639] ^ cw[1641] ^ cw[1643] ^ cw[1645] ^ cw[1647] ^ cw[1649] ^ cw[1651] ^ cw[1653] ^ cw[1655] ^ cw[1657] ^ cw[1659] ^ cw[1661] ^ cw[1663] ^ cw[1665] ^ cw[1667] ^ cw[1669] ^ cw[1671] ^ cw[1673] ^ cw[1675] ^ cw[1677] ^ cw[1679] ^ cw[1681] ^ cw[1683] ^ cw[1685] ^ cw[1687] ^ cw[1689] ^ cw[1691] ^ cw[1693] ^ cw[1695] ^ cw[1697] ^ cw[1699] ^ cw[1701] ^ cw[1703] ^ cw[1705] ^ cw[1707] ^ cw[1709] ^ cw[1711] ^ cw[1713] ^ cw[1715] ^ cw[1717] ^ cw[1719] ^ cw[1721] ^ cw[1723] ^ cw[1725] ^ cw[1727] ^ cw[1729] ^ cw[1731] ^ cw[1733] ^ cw[1735] ^ cw[1737] ^ cw[1739] ^ cw[1741] ^ cw[1743] ^ cw[1745] ^ cw[1747] ^ cw[1749] ^ cw[1751] ^ cw[1753] ^ cw[1755] ^ cw[1757] ^ cw[1759] ^ cw[1761] ^ cw[1763] ^ cw[1765] ^ cw[1767] ^ cw[1769] ^ cw[1771] ^ cw[1773] ^ cw[1775] ^ cw[1777] ^ cw[1779] ^ cw[1781] ^ cw[1783] ^ cw[1785] ^ cw[1787] ^ cw[1789] ^ cw[1791] ^ cw[1793] ^ cw[1795] ^ cw[1797] ^ cw[1799] ^ cw[1801] ^ cw[1803] ^ cw[1805] ^ cw[1807] ^ cw[1809] ^ cw[1811] ^ cw[1813] ^ cw[1815] ^ cw[1817] ^ cw[1819] ^ cw[1821] ^ cw[1823] ^ cw[1825] ^ cw[1827] ^ cw[1829] ^ cw[1831] ^ cw[1833] ^ cw[1835] ^ cw[1837] ^ cw[1839] ^ cw[1841] ^ cw[1843] ^ cw[1845] ^ cw[1847] ^ cw[1849] ^ cw[1851] ^ cw[1853] ^ cw[1855] ^ cw[1857] ^ cw[1859] ^ cw[1861] ^ cw[1863] ^ cw[1865] ^ cw[1867] ^ cw[1869] ^ cw[1871] ^ cw[1873] ^ cw[1875] ^ cw[1877] ^ cw[1879] ^ cw[1881] ^ cw[1883] ^ cw[1885] ^ cw[1887] ^ cw[1889] ^ cw[1891] ^ cw[1893] ^ cw[1895] ^ cw[1897] ^ cw[1899] ^ cw[1901] ^ cw[1903] ^ cw[1905] ^ cw[1907] ^ cw[1909] ^ cw[1911] ^ cw[1913] ^ cw[1915] ^ cw[1917] ^ cw[1919] ^ cw[1921] ^ cw[1923] ^ cw[1925] ^ cw[1927] ^ cw[1929] ^ cw[1931] ^ cw[1933] ^ cw[1935] ^ cw[1937] ^ cw[1939] ^ cw[1941] ^ cw[1943] ^ cw[1945] ^ cw[1947] ^ cw[1949] ^ cw[1951] ^ cw[1953] ^ cw[1955] ^ cw[1957] ^ cw[1959] ^ cw[1961] ^ cw[1963] ^ cw[1965] ^ cw[1967] ^ cw[1969] ^ cw[1971] ^ cw[1973] ^ cw[1975] ^ cw[1977] ^ cw[1979] ^ cw[1981] ^ cw[1983] ^ cw[1985] ^ cw[1987] ^ cw[1989] ^ cw[1991] ^ cw[1993] ^ cw[1995] ^ cw[1997] ^ cw[1999] ^ cw[2001] ^ cw[2003] ^ cw[2005] ^ cw[2007] ^ cw[2009] ^ cw[2011] ^ cw[2013] ^ cw[2015] ^ cw[2017] ^ cw[2019] ^ cw[2021] ^ cw[2023] ^ cw[2024] ^ cw[2025] ^ cw[2026] ^ cw[2027] ^ cw[2028] ^ cw[2029] ^ cw[2030] ^ cw[2031] ^ cw[2032] ^ cw[2033] ^ cw[2034] ^ cw[2047];
    assign parity_check_matrix[0] = 12'b000000000111;
    assign parity_check_matrix[1] = 12'b111111111000;
    assign parity_check_matrix[2] = 12'b000000001011;
    assign parity_check_matrix[3] = 12'b111111110100;
    assign parity_check_matrix[4] = 12'b000000010011;
    assign parity_check_matrix[5] = 12'b111111101100;
    assign parity_check_matrix[6] = 12'b000000100011;
    assign parity_check_matrix[7] = 12'b111111011100;
    assign parity_check_matrix[8] = 12'b000001000011;
    assign parity_check_matrix[9] = 12'b111110111100;
    assign parity_check_matrix[10] = 12'b000010000011;
    assign parity_check_matrix[11] = 12'b111101111100;
    assign parity_check_matrix[12] = 12'b000100000011;
    assign parity_check_matrix[13] = 12'b111011111100;
    assign parity_check_matrix[14] = 12'b001000000011;
    assign parity_check_matrix[15] = 12'b110111111100;
    assign parity_check_matrix[16] = 12'b010000000011;
    assign parity_check_matrix[17] = 12'b101111111100;
    assign parity_check_matrix[18] = 12'b100000000011;
    assign parity_check_matrix[19] = 12'b011111111100;
    assign parity_check_matrix[20] = 12'b000000001101;
    assign parity_check_matrix[21] = 12'b111111110010;
    assign parity_check_matrix[22] = 12'b000000010101;
    assign parity_check_matrix[23] = 12'b111111101010;
    assign parity_check_matrix[24] = 12'b000000100101;
    assign parity_check_matrix[25] = 12'b111111011010;
    assign parity_check_matrix[26] = 12'b000001000101;
    assign parity_check_matrix[27] = 12'b111110111010;
    assign parity_check_matrix[28] = 12'b000010000101;
    assign parity_check_matrix[29] = 12'b111101111010;
    assign parity_check_matrix[30] = 12'b000100000101;
    assign parity_check_matrix[31] = 12'b111011111010;
    assign parity_check_matrix[32] = 12'b001000000101;
    assign parity_check_matrix[33] = 12'b110111111010;
    assign parity_check_matrix[34] = 12'b010000000101;
    assign parity_check_matrix[35] = 12'b101111111010;
    assign parity_check_matrix[36] = 12'b100000000101;
    assign parity_check_matrix[37] = 12'b011111111010;
    assign parity_check_matrix[38] = 12'b000000011001;
    assign parity_check_matrix[39] = 12'b111111100110;
    assign parity_check_matrix[40] = 12'b000000101001;
    assign parity_check_matrix[41] = 12'b111111010110;
    assign parity_check_matrix[42] = 12'b000001001001;
    assign parity_check_matrix[43] = 12'b111110110110;
    assign parity_check_matrix[44] = 12'b000010001001;
    assign parity_check_matrix[45] = 12'b111101110110;
    assign parity_check_matrix[46] = 12'b000100001001;
    assign parity_check_matrix[47] = 12'b111011110110;
    assign parity_check_matrix[48] = 12'b001000001001;
    assign parity_check_matrix[49] = 12'b110111110110;
    assign parity_check_matrix[50] = 12'b010000001001;
    assign parity_check_matrix[51] = 12'b101111110110;
    assign parity_check_matrix[52] = 12'b100000001001;
    assign parity_check_matrix[53] = 12'b011111110110;
    assign parity_check_matrix[54] = 12'b000000110001;
    assign parity_check_matrix[55] = 12'b111111001110;
    assign parity_check_matrix[56] = 12'b000001010001;
    assign parity_check_matrix[57] = 12'b111110101110;
    assign parity_check_matrix[58] = 12'b000010010001;
    assign parity_check_matrix[59] = 12'b111101101110;
    assign parity_check_matrix[60] = 12'b000100010001;
    assign parity_check_matrix[61] = 12'b111011101110;
    assign parity_check_matrix[62] = 12'b001000010001;
    assign parity_check_matrix[63] = 12'b110111101110;
    assign parity_check_matrix[64] = 12'b010000010001;
    assign parity_check_matrix[65] = 12'b101111101110;
    assign parity_check_matrix[66] = 12'b100000010001;
    assign parity_check_matrix[67] = 12'b011111101110;
    assign parity_check_matrix[68] = 12'b000001100001;
    assign parity_check_matrix[69] = 12'b111110011110;
    assign parity_check_matrix[70] = 12'b000010100001;
    assign parity_check_matrix[71] = 12'b111101011110;
    assign parity_check_matrix[72] = 12'b000100100001;
    assign parity_check_matrix[73] = 12'b111011011110;
    assign parity_check_matrix[74] = 12'b001000100001;
    assign parity_check_matrix[75] = 12'b110111011110;
    assign parity_check_matrix[76] = 12'b010000100001;
    assign parity_check_matrix[77] = 12'b101111011110;
    assign parity_check_matrix[78] = 12'b100000100001;
    assign parity_check_matrix[79] = 12'b011111011110;
    assign parity_check_matrix[80] = 12'b000011000001;
    assign parity_check_matrix[81] = 12'b111100111110;
    assign parity_check_matrix[82] = 12'b000101000001;
    assign parity_check_matrix[83] = 12'b111010111110;
    assign parity_check_matrix[84] = 12'b001001000001;
    assign parity_check_matrix[85] = 12'b110110111110;
    assign parity_check_matrix[86] = 12'b010001000001;
    assign parity_check_matrix[87] = 12'b101110111110;
    assign parity_check_matrix[88] = 12'b100001000001;
    assign parity_check_matrix[89] = 12'b011110111110;
    assign parity_check_matrix[90] = 12'b000110000001;
    assign parity_check_matrix[91] = 12'b111001111110;
    assign parity_check_matrix[92] = 12'b001010000001;
    assign parity_check_matrix[93] = 12'b110101111110;
    assign parity_check_matrix[94] = 12'b010010000001;
    assign parity_check_matrix[95] = 12'b101101111110;
    assign parity_check_matrix[96] = 12'b100010000001;
    assign parity_check_matrix[97] = 12'b011101111110;
    assign parity_check_matrix[98] = 12'b001100000001;
    assign parity_check_matrix[99] = 12'b110011111110;
    assign parity_check_matrix[100] = 12'b010100000001;
    assign parity_check_matrix[101] = 12'b101011111110;
    assign parity_check_matrix[102] = 12'b100100000001;
    assign parity_check_matrix[103] = 12'b011011111110;
    assign parity_check_matrix[104] = 12'b011000000001;
    assign parity_check_matrix[105] = 12'b100111111110;
    assign parity_check_matrix[106] = 12'b101000000001;
    assign parity_check_matrix[107] = 12'b010111111110;
    assign parity_check_matrix[108] = 12'b110000000001;
    assign parity_check_matrix[109] = 12'b001111111110;
    assign parity_check_matrix[110] = 12'b000000001110;
    assign parity_check_matrix[111] = 12'b111111110001;
    assign parity_check_matrix[112] = 12'b000000010110;
    assign parity_check_matrix[113] = 12'b111111101001;
    assign parity_check_matrix[114] = 12'b000000100110;
    assign parity_check_matrix[115] = 12'b111111011001;
    assign parity_check_matrix[116] = 12'b000001000110;
    assign parity_check_matrix[117] = 12'b111110111001;
    assign parity_check_matrix[118] = 12'b000010000110;
    assign parity_check_matrix[119] = 12'b111101111001;
    assign parity_check_matrix[120] = 12'b000100000110;
    assign parity_check_matrix[121] = 12'b111011111001;
    assign parity_check_matrix[122] = 12'b001000000110;
    assign parity_check_matrix[123] = 12'b110111111001;
    assign parity_check_matrix[124] = 12'b010000000110;
    assign parity_check_matrix[125] = 12'b101111111001;
    assign parity_check_matrix[126] = 12'b100000000110;
    assign parity_check_matrix[127] = 12'b011111111001;
    assign parity_check_matrix[128] = 12'b000000011010;
    assign parity_check_matrix[129] = 12'b111111100101;
    assign parity_check_matrix[130] = 12'b000000101010;
    assign parity_check_matrix[131] = 12'b111111010101;
    assign parity_check_matrix[132] = 12'b000001001010;
    assign parity_check_matrix[133] = 12'b111110110101;
    assign parity_check_matrix[134] = 12'b000010001010;
    assign parity_check_matrix[135] = 12'b111101110101;
    assign parity_check_matrix[136] = 12'b000100001010;
    assign parity_check_matrix[137] = 12'b111011110101;
    assign parity_check_matrix[138] = 12'b001000001010;
    assign parity_check_matrix[139] = 12'b110111110101;
    assign parity_check_matrix[140] = 12'b010000001010;
    assign parity_check_matrix[141] = 12'b101111110101;
    assign parity_check_matrix[142] = 12'b100000001010;
    assign parity_check_matrix[143] = 12'b011111110101;
    assign parity_check_matrix[144] = 12'b000000110010;
    assign parity_check_matrix[145] = 12'b111111001101;
    assign parity_check_matrix[146] = 12'b000001010010;
    assign parity_check_matrix[147] = 12'b111110101101;
    assign parity_check_matrix[148] = 12'b000010010010;
    assign parity_check_matrix[149] = 12'b111101101101;
    assign parity_check_matrix[150] = 12'b000100010010;
    assign parity_check_matrix[151] = 12'b111011101101;
    assign parity_check_matrix[152] = 12'b001000010010;
    assign parity_check_matrix[153] = 12'b110111101101;
    assign parity_check_matrix[154] = 12'b010000010010;
    assign parity_check_matrix[155] = 12'b101111101101;
    assign parity_check_matrix[156] = 12'b100000010010;
    assign parity_check_matrix[157] = 12'b011111101101;
    assign parity_check_matrix[158] = 12'b000001100010;
    assign parity_check_matrix[159] = 12'b111110011101;
    assign parity_check_matrix[160] = 12'b000010100010;
    assign parity_check_matrix[161] = 12'b111101011101;
    assign parity_check_matrix[162] = 12'b000100100010;
    assign parity_check_matrix[163] = 12'b111011011101;
    assign parity_check_matrix[164] = 12'b001000100010;
    assign parity_check_matrix[165] = 12'b110111011101;
    assign parity_check_matrix[166] = 12'b010000100010;
    assign parity_check_matrix[167] = 12'b101111011101;
    assign parity_check_matrix[168] = 12'b100000100010;
    assign parity_check_matrix[169] = 12'b011111011101;
    assign parity_check_matrix[170] = 12'b000011000010;
    assign parity_check_matrix[171] = 12'b111100111101;
    assign parity_check_matrix[172] = 12'b000101000010;
    assign parity_check_matrix[173] = 12'b111010111101;
    assign parity_check_matrix[174] = 12'b001001000010;
    assign parity_check_matrix[175] = 12'b110110111101;
    assign parity_check_matrix[176] = 12'b010001000010;
    assign parity_check_matrix[177] = 12'b101110111101;
    assign parity_check_matrix[178] = 12'b100001000010;
    assign parity_check_matrix[179] = 12'b011110111101;
    assign parity_check_matrix[180] = 12'b000110000010;
    assign parity_check_matrix[181] = 12'b111001111101;
    assign parity_check_matrix[182] = 12'b001010000010;
    assign parity_check_matrix[183] = 12'b110101111101;
    assign parity_check_matrix[184] = 12'b010010000010;
    assign parity_check_matrix[185] = 12'b101101111101;
    assign parity_check_matrix[186] = 12'b100010000010;
    assign parity_check_matrix[187] = 12'b011101111101;
    assign parity_check_matrix[188] = 12'b001100000010;
    assign parity_check_matrix[189] = 12'b110011111101;
    assign parity_check_matrix[190] = 12'b010100000010;
    assign parity_check_matrix[191] = 12'b101011111101;
    assign parity_check_matrix[192] = 12'b100100000010;
    assign parity_check_matrix[193] = 12'b011011111101;
    assign parity_check_matrix[194] = 12'b011000000010;
    assign parity_check_matrix[195] = 12'b100111111101;
    assign parity_check_matrix[196] = 12'b101000000010;
    assign parity_check_matrix[197] = 12'b010111111101;
    assign parity_check_matrix[198] = 12'b110000000010;
    assign parity_check_matrix[199] = 12'b001111111101;
    assign parity_check_matrix[200] = 12'b000000011100;
    assign parity_check_matrix[201] = 12'b111111100011;
    assign parity_check_matrix[202] = 12'b000000101100;
    assign parity_check_matrix[203] = 12'b111111010011;
    assign parity_check_matrix[204] = 12'b000001001100;
    assign parity_check_matrix[205] = 12'b111110110011;
    assign parity_check_matrix[206] = 12'b000010001100;
    assign parity_check_matrix[207] = 12'b111101110011;
    assign parity_check_matrix[208] = 12'b000100001100;
    assign parity_check_matrix[209] = 12'b111011110011;
    assign parity_check_matrix[210] = 12'b001000001100;
    assign parity_check_matrix[211] = 12'b110111110011;
    assign parity_check_matrix[212] = 12'b010000001100;
    assign parity_check_matrix[213] = 12'b101111110011;
    assign parity_check_matrix[214] = 12'b100000001100;
    assign parity_check_matrix[215] = 12'b011111110011;
    assign parity_check_matrix[216] = 12'b000000110100;
    assign parity_check_matrix[217] = 12'b111111001011;
    assign parity_check_matrix[218] = 12'b000001010100;
    assign parity_check_matrix[219] = 12'b111110101011;
    assign parity_check_matrix[220] = 12'b000010010100;
    assign parity_check_matrix[221] = 12'b111101101011;
    assign parity_check_matrix[222] = 12'b000100010100;
    assign parity_check_matrix[223] = 12'b111011101011;
    assign parity_check_matrix[224] = 12'b001000010100;
    assign parity_check_matrix[225] = 12'b110111101011;
    assign parity_check_matrix[226] = 12'b010000010100;
    assign parity_check_matrix[227] = 12'b101111101011;
    assign parity_check_matrix[228] = 12'b100000010100;
    assign parity_check_matrix[229] = 12'b011111101011;
    assign parity_check_matrix[230] = 12'b000001100100;
    assign parity_check_matrix[231] = 12'b111110011011;
    assign parity_check_matrix[232] = 12'b000010100100;
    assign parity_check_matrix[233] = 12'b111101011011;
    assign parity_check_matrix[234] = 12'b000100100100;
    assign parity_check_matrix[235] = 12'b111011011011;
    assign parity_check_matrix[236] = 12'b001000100100;
    assign parity_check_matrix[237] = 12'b110111011011;
    assign parity_check_matrix[238] = 12'b010000100100;
    assign parity_check_matrix[239] = 12'b101111011011;
    assign parity_check_matrix[240] = 12'b100000100100;
    assign parity_check_matrix[241] = 12'b011111011011;
    assign parity_check_matrix[242] = 12'b000011000100;
    assign parity_check_matrix[243] = 12'b111100111011;
    assign parity_check_matrix[244] = 12'b000101000100;
    assign parity_check_matrix[245] = 12'b111010111011;
    assign parity_check_matrix[246] = 12'b001001000100;
    assign parity_check_matrix[247] = 12'b110110111011;
    assign parity_check_matrix[248] = 12'b010001000100;
    assign parity_check_matrix[249] = 12'b101110111011;
    assign parity_check_matrix[250] = 12'b100001000100;
    assign parity_check_matrix[251] = 12'b011110111011;
    assign parity_check_matrix[252] = 12'b000110000100;
    assign parity_check_matrix[253] = 12'b111001111011;
    assign parity_check_matrix[254] = 12'b001010000100;
    assign parity_check_matrix[255] = 12'b110101111011;
    assign parity_check_matrix[256] = 12'b010010000100;
    assign parity_check_matrix[257] = 12'b101101111011;
    assign parity_check_matrix[258] = 12'b100010000100;
    assign parity_check_matrix[259] = 12'b011101111011;
    assign parity_check_matrix[260] = 12'b001100000100;
    assign parity_check_matrix[261] = 12'b110011111011;
    assign parity_check_matrix[262] = 12'b010100000100;
    assign parity_check_matrix[263] = 12'b101011111011;
    assign parity_check_matrix[264] = 12'b100100000100;
    assign parity_check_matrix[265] = 12'b011011111011;
    assign parity_check_matrix[266] = 12'b011000000100;
    assign parity_check_matrix[267] = 12'b100111111011;
    assign parity_check_matrix[268] = 12'b101000000100;
    assign parity_check_matrix[269] = 12'b010111111011;
    assign parity_check_matrix[270] = 12'b110000000100;
    assign parity_check_matrix[271] = 12'b001111111011;
    assign parity_check_matrix[272] = 12'b000000111000;
    assign parity_check_matrix[273] = 12'b111111000111;
    assign parity_check_matrix[274] = 12'b000001011000;
    assign parity_check_matrix[275] = 12'b111110100111;
    assign parity_check_matrix[276] = 12'b000010011000;
    assign parity_check_matrix[277] = 12'b111101100111;
    assign parity_check_matrix[278] = 12'b000100011000;
    assign parity_check_matrix[279] = 12'b111011100111;
    assign parity_check_matrix[280] = 12'b001000011000;
    assign parity_check_matrix[281] = 12'b110111100111;
    assign parity_check_matrix[282] = 12'b010000011000;
    assign parity_check_matrix[283] = 12'b101111100111;
    assign parity_check_matrix[284] = 12'b100000011000;
    assign parity_check_matrix[285] = 12'b011111100111;
    assign parity_check_matrix[286] = 12'b000001101000;
    assign parity_check_matrix[287] = 12'b111110010111;
    assign parity_check_matrix[288] = 12'b000010101000;
    assign parity_check_matrix[289] = 12'b111101010111;
    assign parity_check_matrix[290] = 12'b000100101000;
    assign parity_check_matrix[291] = 12'b111011010111;
    assign parity_check_matrix[292] = 12'b001000101000;
    assign parity_check_matrix[293] = 12'b110111010111;
    assign parity_check_matrix[294] = 12'b010000101000;
    assign parity_check_matrix[295] = 12'b101111010111;
    assign parity_check_matrix[296] = 12'b100000101000;
    assign parity_check_matrix[297] = 12'b011111010111;
    assign parity_check_matrix[298] = 12'b000011001000;
    assign parity_check_matrix[299] = 12'b111100110111;
    assign parity_check_matrix[300] = 12'b000101001000;
    assign parity_check_matrix[301] = 12'b111010110111;
    assign parity_check_matrix[302] = 12'b001001001000;
    assign parity_check_matrix[303] = 12'b110110110111;
    assign parity_check_matrix[304] = 12'b010001001000;
    assign parity_check_matrix[305] = 12'b101110110111;
    assign parity_check_matrix[306] = 12'b100001001000;
    assign parity_check_matrix[307] = 12'b011110110111;
    assign parity_check_matrix[308] = 12'b000110001000;
    assign parity_check_matrix[309] = 12'b111001110111;
    assign parity_check_matrix[310] = 12'b001010001000;
    assign parity_check_matrix[311] = 12'b110101110111;
    assign parity_check_matrix[312] = 12'b010010001000;
    assign parity_check_matrix[313] = 12'b101101110111;
    assign parity_check_matrix[314] = 12'b100010001000;
    assign parity_check_matrix[315] = 12'b011101110111;
    assign parity_check_matrix[316] = 12'b001100001000;
    assign parity_check_matrix[317] = 12'b110011110111;
    assign parity_check_matrix[318] = 12'b010100001000;
    assign parity_check_matrix[319] = 12'b101011110111;
    assign parity_check_matrix[320] = 12'b100100001000;
    assign parity_check_matrix[321] = 12'b011011110111;
    assign parity_check_matrix[322] = 12'b011000001000;
    assign parity_check_matrix[323] = 12'b100111110111;
    assign parity_check_matrix[324] = 12'b101000001000;
    assign parity_check_matrix[325] = 12'b010111110111;
    assign parity_check_matrix[326] = 12'b110000001000;
    assign parity_check_matrix[327] = 12'b001111110111;
    assign parity_check_matrix[328] = 12'b000001110000;
    assign parity_check_matrix[329] = 12'b111110001111;
    assign parity_check_matrix[330] = 12'b000010110000;
    assign parity_check_matrix[331] = 12'b111101001111;
    assign parity_check_matrix[332] = 12'b000100110000;
    assign parity_check_matrix[333] = 12'b111011001111;
    assign parity_check_matrix[334] = 12'b001000110000;
    assign parity_check_matrix[335] = 12'b110111001111;
    assign parity_check_matrix[336] = 12'b010000110000;
    assign parity_check_matrix[337] = 12'b101111001111;
    assign parity_check_matrix[338] = 12'b100000110000;
    assign parity_check_matrix[339] = 12'b011111001111;
    assign parity_check_matrix[340] = 12'b000011010000;
    assign parity_check_matrix[341] = 12'b111100101111;
    assign parity_check_matrix[342] = 12'b000101010000;
    assign parity_check_matrix[343] = 12'b111010101111;
    assign parity_check_matrix[344] = 12'b001001010000;
    assign parity_check_matrix[345] = 12'b110110101111;
    assign parity_check_matrix[346] = 12'b010001010000;
    assign parity_check_matrix[347] = 12'b101110101111;
    assign parity_check_matrix[348] = 12'b100001010000;
    assign parity_check_matrix[349] = 12'b011110101111;
    assign parity_check_matrix[350] = 12'b000110010000;
    assign parity_check_matrix[351] = 12'b111001101111;
    assign parity_check_matrix[352] = 12'b001010010000;
    assign parity_check_matrix[353] = 12'b110101101111;
    assign parity_check_matrix[354] = 12'b010010010000;
    assign parity_check_matrix[355] = 12'b101101101111;
    assign parity_check_matrix[356] = 12'b100010010000;
    assign parity_check_matrix[357] = 12'b011101101111;
    assign parity_check_matrix[358] = 12'b001100010000;
    assign parity_check_matrix[359] = 12'b110011101111;
    assign parity_check_matrix[360] = 12'b010100010000;
    assign parity_check_matrix[361] = 12'b101011101111;
    assign parity_check_matrix[362] = 12'b100100010000;
    assign parity_check_matrix[363] = 12'b011011101111;
    assign parity_check_matrix[364] = 12'b011000010000;
    assign parity_check_matrix[365] = 12'b100111101111;
    assign parity_check_matrix[366] = 12'b101000010000;
    assign parity_check_matrix[367] = 12'b010111101111;
    assign parity_check_matrix[368] = 12'b110000010000;
    assign parity_check_matrix[369] = 12'b001111101111;
    assign parity_check_matrix[370] = 12'b000011100000;
    assign parity_check_matrix[371] = 12'b111100011111;
    assign parity_check_matrix[372] = 12'b000101100000;
    assign parity_check_matrix[373] = 12'b111010011111;
    assign parity_check_matrix[374] = 12'b001001100000;
    assign parity_check_matrix[375] = 12'b110110011111;
    assign parity_check_matrix[376] = 12'b010001100000;
    assign parity_check_matrix[377] = 12'b101110011111;
    assign parity_check_matrix[378] = 12'b100001100000;
    assign parity_check_matrix[379] = 12'b011110011111;
    assign parity_check_matrix[380] = 12'b000110100000;
    assign parity_check_matrix[381] = 12'b111001011111;
    assign parity_check_matrix[382] = 12'b001010100000;
    assign parity_check_matrix[383] = 12'b110101011111;
    assign parity_check_matrix[384] = 12'b010010100000;
    assign parity_check_matrix[385] = 12'b101101011111;
    assign parity_check_matrix[386] = 12'b100010100000;
    assign parity_check_matrix[387] = 12'b011101011111;
    assign parity_check_matrix[388] = 12'b001100100000;
    assign parity_check_matrix[389] = 12'b110011011111;
    assign parity_check_matrix[390] = 12'b010100100000;
    assign parity_check_matrix[391] = 12'b101011011111;
    assign parity_check_matrix[392] = 12'b100100100000;
    assign parity_check_matrix[393] = 12'b011011011111;
    assign parity_check_matrix[394] = 12'b011000100000;
    assign parity_check_matrix[395] = 12'b100111011111;
    assign parity_check_matrix[396] = 12'b101000100000;
    assign parity_check_matrix[397] = 12'b010111011111;
    assign parity_check_matrix[398] = 12'b110000100000;
    assign parity_check_matrix[399] = 12'b001111011111;
    assign parity_check_matrix[400] = 12'b000111000000;
    assign parity_check_matrix[401] = 12'b111000111111;
    assign parity_check_matrix[402] = 12'b001011000000;
    assign parity_check_matrix[403] = 12'b110100111111;
    assign parity_check_matrix[404] = 12'b010011000000;
    assign parity_check_matrix[405] = 12'b101100111111;
    assign parity_check_matrix[406] = 12'b100011000000;
    assign parity_check_matrix[407] = 12'b011100111111;
    assign parity_check_matrix[408] = 12'b001101000000;
    assign parity_check_matrix[409] = 12'b110010111111;
    assign parity_check_matrix[410] = 12'b010101000000;
    assign parity_check_matrix[411] = 12'b101010111111;
    assign parity_check_matrix[412] = 12'b100101000000;
    assign parity_check_matrix[413] = 12'b011010111111;
    assign parity_check_matrix[414] = 12'b011001000000;
    assign parity_check_matrix[415] = 12'b100110111111;
    assign parity_check_matrix[416] = 12'b101001000000;
    assign parity_check_matrix[417] = 12'b010110111111;
    assign parity_check_matrix[418] = 12'b110001000000;
    assign parity_check_matrix[419] = 12'b001110111111;
    assign parity_check_matrix[420] = 12'b001110000000;
    assign parity_check_matrix[421] = 12'b110001111111;
    assign parity_check_matrix[422] = 12'b010110000000;
    assign parity_check_matrix[423] = 12'b101001111111;
    assign parity_check_matrix[424] = 12'b100110000000;
    assign parity_check_matrix[425] = 12'b011001111111;
    assign parity_check_matrix[426] = 12'b011010000000;
    assign parity_check_matrix[427] = 12'b100101111111;
    assign parity_check_matrix[428] = 12'b101010000000;
    assign parity_check_matrix[429] = 12'b010101111111;
    assign parity_check_matrix[430] = 12'b110010000000;
    assign parity_check_matrix[431] = 12'b001101111111;
    assign parity_check_matrix[432] = 12'b011100000000;
    assign parity_check_matrix[433] = 12'b100011111111;
    assign parity_check_matrix[434] = 12'b101100000000;
    assign parity_check_matrix[435] = 12'b010011111111;
    assign parity_check_matrix[436] = 12'b110100000000;
    assign parity_check_matrix[437] = 12'b001011111111;
    assign parity_check_matrix[438] = 12'b111000000000;
    assign parity_check_matrix[439] = 12'b000111111111;
    assign parity_check_matrix[440] = 12'b000000011111;
    assign parity_check_matrix[441] = 12'b111111100000;
    assign parity_check_matrix[442] = 12'b000000101111;
    assign parity_check_matrix[443] = 12'b111111010000;
    assign parity_check_matrix[444] = 12'b000001001111;
    assign parity_check_matrix[445] = 12'b111110110000;
    assign parity_check_matrix[446] = 12'b000010001111;
    assign parity_check_matrix[447] = 12'b111101110000;
    assign parity_check_matrix[448] = 12'b000100001111;
    assign parity_check_matrix[449] = 12'b111011110000;
    assign parity_check_matrix[450] = 12'b001000001111;
    assign parity_check_matrix[451] = 12'b110111110000;
    assign parity_check_matrix[452] = 12'b010000001111;
    assign parity_check_matrix[453] = 12'b101111110000;
    assign parity_check_matrix[454] = 12'b100000001111;
    assign parity_check_matrix[455] = 12'b011111110000;
    assign parity_check_matrix[456] = 12'b000000110111;
    assign parity_check_matrix[457] = 12'b111111001000;
    assign parity_check_matrix[458] = 12'b000001010111;
    assign parity_check_matrix[459] = 12'b111110101000;
    assign parity_check_matrix[460] = 12'b000010010111;
    assign parity_check_matrix[461] = 12'b111101101000;
    assign parity_check_matrix[462] = 12'b000100010111;
    assign parity_check_matrix[463] = 12'b111011101000;
    assign parity_check_matrix[464] = 12'b001000010111;
    assign parity_check_matrix[465] = 12'b110111101000;
    assign parity_check_matrix[466] = 12'b010000010111;
    assign parity_check_matrix[467] = 12'b101111101000;
    assign parity_check_matrix[468] = 12'b100000010111;
    assign parity_check_matrix[469] = 12'b011111101000;
    assign parity_check_matrix[470] = 12'b000001100111;
    assign parity_check_matrix[471] = 12'b111110011000;
    assign parity_check_matrix[472] = 12'b000010100111;
    assign parity_check_matrix[473] = 12'b111101011000;
    assign parity_check_matrix[474] = 12'b000100100111;
    assign parity_check_matrix[475] = 12'b111011011000;
    assign parity_check_matrix[476] = 12'b001000100111;
    assign parity_check_matrix[477] = 12'b110111011000;
    assign parity_check_matrix[478] = 12'b010000100111;
    assign parity_check_matrix[479] = 12'b101111011000;
    assign parity_check_matrix[480] = 12'b100000100111;
    assign parity_check_matrix[481] = 12'b011111011000;
    assign parity_check_matrix[482] = 12'b000011000111;
    assign parity_check_matrix[483] = 12'b111100111000;
    assign parity_check_matrix[484] = 12'b000101000111;
    assign parity_check_matrix[485] = 12'b111010111000;
    assign parity_check_matrix[486] = 12'b001001000111;
    assign parity_check_matrix[487] = 12'b110110111000;
    assign parity_check_matrix[488] = 12'b010001000111;
    assign parity_check_matrix[489] = 12'b101110111000;
    assign parity_check_matrix[490] = 12'b100001000111;
    assign parity_check_matrix[491] = 12'b011110111000;
    assign parity_check_matrix[492] = 12'b000110000111;
    assign parity_check_matrix[493] = 12'b111001111000;
    assign parity_check_matrix[494] = 12'b001010000111;
    assign parity_check_matrix[495] = 12'b110101111000;
    assign parity_check_matrix[496] = 12'b010010000111;
    assign parity_check_matrix[497] = 12'b101101111000;
    assign parity_check_matrix[498] = 12'b100010000111;
    assign parity_check_matrix[499] = 12'b011101111000;
    assign parity_check_matrix[500] = 12'b001100000111;
    assign parity_check_matrix[501] = 12'b110011111000;
    assign parity_check_matrix[502] = 12'b010100000111;
    assign parity_check_matrix[503] = 12'b101011111000;
    assign parity_check_matrix[504] = 12'b100100000111;
    assign parity_check_matrix[505] = 12'b011011111000;
    assign parity_check_matrix[506] = 12'b011000000111;
    assign parity_check_matrix[507] = 12'b100111111000;
    assign parity_check_matrix[508] = 12'b101000000111;
    assign parity_check_matrix[509] = 12'b010111111000;
    assign parity_check_matrix[510] = 12'b110000000111;
    assign parity_check_matrix[511] = 12'b001111111000;
    assign parity_check_matrix[512] = 12'b000000111011;
    assign parity_check_matrix[513] = 12'b111111000100;
    assign parity_check_matrix[514] = 12'b000001011011;
    assign parity_check_matrix[515] = 12'b111110100100;
    assign parity_check_matrix[516] = 12'b000010011011;
    assign parity_check_matrix[517] = 12'b111101100100;
    assign parity_check_matrix[518] = 12'b000100011011;
    assign parity_check_matrix[519] = 12'b111011100100;
    assign parity_check_matrix[520] = 12'b001000011011;
    assign parity_check_matrix[521] = 12'b110111100100;
    assign parity_check_matrix[522] = 12'b010000011011;
    assign parity_check_matrix[523] = 12'b101111100100;
    assign parity_check_matrix[524] = 12'b100000011011;
    assign parity_check_matrix[525] = 12'b011111100100;
    assign parity_check_matrix[526] = 12'b000001101011;
    assign parity_check_matrix[527] = 12'b111110010100;
    assign parity_check_matrix[528] = 12'b000010101011;
    assign parity_check_matrix[529] = 12'b111101010100;
    assign parity_check_matrix[530] = 12'b000100101011;
    assign parity_check_matrix[531] = 12'b111011010100;
    assign parity_check_matrix[532] = 12'b001000101011;
    assign parity_check_matrix[533] = 12'b110111010100;
    assign parity_check_matrix[534] = 12'b010000101011;
    assign parity_check_matrix[535] = 12'b101111010100;
    assign parity_check_matrix[536] = 12'b100000101011;
    assign parity_check_matrix[537] = 12'b011111010100;
    assign parity_check_matrix[538] = 12'b000011001011;
    assign parity_check_matrix[539] = 12'b111100110100;
    assign parity_check_matrix[540] = 12'b000101001011;
    assign parity_check_matrix[541] = 12'b111010110100;
    assign parity_check_matrix[542] = 12'b001001001011;
    assign parity_check_matrix[543] = 12'b110110110100;
    assign parity_check_matrix[544] = 12'b010001001011;
    assign parity_check_matrix[545] = 12'b101110110100;
    assign parity_check_matrix[546] = 12'b100001001011;
    assign parity_check_matrix[547] = 12'b011110110100;
    assign parity_check_matrix[548] = 12'b000110001011;
    assign parity_check_matrix[549] = 12'b111001110100;
    assign parity_check_matrix[550] = 12'b001010001011;
    assign parity_check_matrix[551] = 12'b110101110100;
    assign parity_check_matrix[552] = 12'b010010001011;
    assign parity_check_matrix[553] = 12'b101101110100;
    assign parity_check_matrix[554] = 12'b100010001011;
    assign parity_check_matrix[555] = 12'b011101110100;
    assign parity_check_matrix[556] = 12'b001100001011;
    assign parity_check_matrix[557] = 12'b110011110100;
    assign parity_check_matrix[558] = 12'b010100001011;
    assign parity_check_matrix[559] = 12'b101011110100;
    assign parity_check_matrix[560] = 12'b100100001011;
    assign parity_check_matrix[561] = 12'b011011110100;
    assign parity_check_matrix[562] = 12'b011000001011;
    assign parity_check_matrix[563] = 12'b100111110100;
    assign parity_check_matrix[564] = 12'b101000001011;
    assign parity_check_matrix[565] = 12'b010111110100;
    assign parity_check_matrix[566] = 12'b110000001011;
    assign parity_check_matrix[567] = 12'b001111110100;
    assign parity_check_matrix[568] = 12'b000001110011;
    assign parity_check_matrix[569] = 12'b111110001100;
    assign parity_check_matrix[570] = 12'b000010110011;
    assign parity_check_matrix[571] = 12'b111101001100;
    assign parity_check_matrix[572] = 12'b000100110011;
    assign parity_check_matrix[573] = 12'b111011001100;
    assign parity_check_matrix[574] = 12'b001000110011;
    assign parity_check_matrix[575] = 12'b110111001100;
    assign parity_check_matrix[576] = 12'b010000110011;
    assign parity_check_matrix[577] = 12'b101111001100;
    assign parity_check_matrix[578] = 12'b100000110011;
    assign parity_check_matrix[579] = 12'b011111001100;
    assign parity_check_matrix[580] = 12'b000011010011;
    assign parity_check_matrix[581] = 12'b111100101100;
    assign parity_check_matrix[582] = 12'b000101010011;
    assign parity_check_matrix[583] = 12'b111010101100;
    assign parity_check_matrix[584] = 12'b001001010011;
    assign parity_check_matrix[585] = 12'b110110101100;
    assign parity_check_matrix[586] = 12'b010001010011;
    assign parity_check_matrix[587] = 12'b101110101100;
    assign parity_check_matrix[588] = 12'b100001010011;
    assign parity_check_matrix[589] = 12'b011110101100;
    assign parity_check_matrix[590] = 12'b000110010011;
    assign parity_check_matrix[591] = 12'b111001101100;
    assign parity_check_matrix[592] = 12'b001010010011;
    assign parity_check_matrix[593] = 12'b110101101100;
    assign parity_check_matrix[594] = 12'b010010010011;
    assign parity_check_matrix[595] = 12'b101101101100;
    assign parity_check_matrix[596] = 12'b100010010011;
    assign parity_check_matrix[597] = 12'b011101101100;
    assign parity_check_matrix[598] = 12'b001100010011;
    assign parity_check_matrix[599] = 12'b110011101100;
    assign parity_check_matrix[600] = 12'b010100010011;
    assign parity_check_matrix[601] = 12'b101011101100;
    assign parity_check_matrix[602] = 12'b100100010011;
    assign parity_check_matrix[603] = 12'b011011101100;
    assign parity_check_matrix[604] = 12'b011000010011;
    assign parity_check_matrix[605] = 12'b100111101100;
    assign parity_check_matrix[606] = 12'b101000010011;
    assign parity_check_matrix[607] = 12'b010111101100;
    assign parity_check_matrix[608] = 12'b110000010011;
    assign parity_check_matrix[609] = 12'b001111101100;
    assign parity_check_matrix[610] = 12'b000011100011;
    assign parity_check_matrix[611] = 12'b111100011100;
    assign parity_check_matrix[612] = 12'b000101100011;
    assign parity_check_matrix[613] = 12'b111010011100;
    assign parity_check_matrix[614] = 12'b001001100011;
    assign parity_check_matrix[615] = 12'b110110011100;
    assign parity_check_matrix[616] = 12'b010001100011;
    assign parity_check_matrix[617] = 12'b101110011100;
    assign parity_check_matrix[618] = 12'b100001100011;
    assign parity_check_matrix[619] = 12'b011110011100;
    assign parity_check_matrix[620] = 12'b000110100011;
    assign parity_check_matrix[621] = 12'b111001011100;
    assign parity_check_matrix[622] = 12'b001010100011;
    assign parity_check_matrix[623] = 12'b110101011100;
    assign parity_check_matrix[624] = 12'b010010100011;
    assign parity_check_matrix[625] = 12'b101101011100;
    assign parity_check_matrix[626] = 12'b100010100011;
    assign parity_check_matrix[627] = 12'b011101011100;
    assign parity_check_matrix[628] = 12'b001100100011;
    assign parity_check_matrix[629] = 12'b110011011100;
    assign parity_check_matrix[630] = 12'b010100100011;
    assign parity_check_matrix[631] = 12'b101011011100;
    assign parity_check_matrix[632] = 12'b100100100011;
    assign parity_check_matrix[633] = 12'b011011011100;
    assign parity_check_matrix[634] = 12'b011000100011;
    assign parity_check_matrix[635] = 12'b100111011100;
    assign parity_check_matrix[636] = 12'b101000100011;
    assign parity_check_matrix[637] = 12'b010111011100;
    assign parity_check_matrix[638] = 12'b110000100011;
    assign parity_check_matrix[639] = 12'b001111011100;
    assign parity_check_matrix[640] = 12'b000111000011;
    assign parity_check_matrix[641] = 12'b111000111100;
    assign parity_check_matrix[642] = 12'b001011000011;
    assign parity_check_matrix[643] = 12'b110100111100;
    assign parity_check_matrix[644] = 12'b010011000011;
    assign parity_check_matrix[645] = 12'b101100111100;
    assign parity_check_matrix[646] = 12'b100011000011;
    assign parity_check_matrix[647] = 12'b011100111100;
    assign parity_check_matrix[648] = 12'b001101000011;
    assign parity_check_matrix[649] = 12'b110010111100;
    assign parity_check_matrix[650] = 12'b010101000011;
    assign parity_check_matrix[651] = 12'b101010111100;
    assign parity_check_matrix[652] = 12'b100101000011;
    assign parity_check_matrix[653] = 12'b011010111100;
    assign parity_check_matrix[654] = 12'b011001000011;
    assign parity_check_matrix[655] = 12'b100110111100;
    assign parity_check_matrix[656] = 12'b101001000011;
    assign parity_check_matrix[657] = 12'b010110111100;
    assign parity_check_matrix[658] = 12'b110001000011;
    assign parity_check_matrix[659] = 12'b001110111100;
    assign parity_check_matrix[660] = 12'b001110000011;
    assign parity_check_matrix[661] = 12'b110001111100;
    assign parity_check_matrix[662] = 12'b010110000011;
    assign parity_check_matrix[663] = 12'b101001111100;
    assign parity_check_matrix[664] = 12'b100110000011;
    assign parity_check_matrix[665] = 12'b011001111100;
    assign parity_check_matrix[666] = 12'b011010000011;
    assign parity_check_matrix[667] = 12'b100101111100;
    assign parity_check_matrix[668] = 12'b101010000011;
    assign parity_check_matrix[669] = 12'b010101111100;
    assign parity_check_matrix[670] = 12'b110010000011;
    assign parity_check_matrix[671] = 12'b001101111100;
    assign parity_check_matrix[672] = 12'b011100000011;
    assign parity_check_matrix[673] = 12'b100011111100;
    assign parity_check_matrix[674] = 12'b101100000011;
    assign parity_check_matrix[675] = 12'b010011111100;
    assign parity_check_matrix[676] = 12'b110100000011;
    assign parity_check_matrix[677] = 12'b001011111100;
    assign parity_check_matrix[678] = 12'b111000000011;
    assign parity_check_matrix[679] = 12'b000111111100;
    assign parity_check_matrix[680] = 12'b000000111101;
    assign parity_check_matrix[681] = 12'b111111000010;
    assign parity_check_matrix[682] = 12'b000001011101;
    assign parity_check_matrix[683] = 12'b111110100010;
    assign parity_check_matrix[684] = 12'b000010011101;
    assign parity_check_matrix[685] = 12'b111101100010;
    assign parity_check_matrix[686] = 12'b000100011101;
    assign parity_check_matrix[687] = 12'b111011100010;
    assign parity_check_matrix[688] = 12'b001000011101;
    assign parity_check_matrix[689] = 12'b110111100010;
    assign parity_check_matrix[690] = 12'b010000011101;
    assign parity_check_matrix[691] = 12'b101111100010;
    assign parity_check_matrix[692] = 12'b100000011101;
    assign parity_check_matrix[693] = 12'b011111100010;
    assign parity_check_matrix[694] = 12'b000001101101;
    assign parity_check_matrix[695] = 12'b111110010010;
    assign parity_check_matrix[696] = 12'b000010101101;
    assign parity_check_matrix[697] = 12'b111101010010;
    assign parity_check_matrix[698] = 12'b000100101101;
    assign parity_check_matrix[699] = 12'b111011010010;
    assign parity_check_matrix[700] = 12'b001000101101;
    assign parity_check_matrix[701] = 12'b110111010010;
    assign parity_check_matrix[702] = 12'b010000101101;
    assign parity_check_matrix[703] = 12'b101111010010;
    assign parity_check_matrix[704] = 12'b100000101101;
    assign parity_check_matrix[705] = 12'b011111010010;
    assign parity_check_matrix[706] = 12'b000011001101;
    assign parity_check_matrix[707] = 12'b111100110010;
    assign parity_check_matrix[708] = 12'b000101001101;
    assign parity_check_matrix[709] = 12'b111010110010;
    assign parity_check_matrix[710] = 12'b001001001101;
    assign parity_check_matrix[711] = 12'b110110110010;
    assign parity_check_matrix[712] = 12'b010001001101;
    assign parity_check_matrix[713] = 12'b101110110010;
    assign parity_check_matrix[714] = 12'b100001001101;
    assign parity_check_matrix[715] = 12'b011110110010;
    assign parity_check_matrix[716] = 12'b000110001101;
    assign parity_check_matrix[717] = 12'b111001110010;
    assign parity_check_matrix[718] = 12'b001010001101;
    assign parity_check_matrix[719] = 12'b110101110010;
    assign parity_check_matrix[720] = 12'b010010001101;
    assign parity_check_matrix[721] = 12'b101101110010;
    assign parity_check_matrix[722] = 12'b100010001101;
    assign parity_check_matrix[723] = 12'b011101110010;
    assign parity_check_matrix[724] = 12'b001100001101;
    assign parity_check_matrix[725] = 12'b110011110010;
    assign parity_check_matrix[726] = 12'b010100001101;
    assign parity_check_matrix[727] = 12'b101011110010;
    assign parity_check_matrix[728] = 12'b100100001101;
    assign parity_check_matrix[729] = 12'b011011110010;
    assign parity_check_matrix[730] = 12'b011000001101;
    assign parity_check_matrix[731] = 12'b100111110010;
    assign parity_check_matrix[732] = 12'b101000001101;
    assign parity_check_matrix[733] = 12'b010111110010;
    assign parity_check_matrix[734] = 12'b110000001101;
    assign parity_check_matrix[735] = 12'b001111110010;
    assign parity_check_matrix[736] = 12'b000001110101;
    assign parity_check_matrix[737] = 12'b111110001010;
    assign parity_check_matrix[738] = 12'b000010110101;
    assign parity_check_matrix[739] = 12'b111101001010;
    assign parity_check_matrix[740] = 12'b000100110101;
    assign parity_check_matrix[741] = 12'b111011001010;
    assign parity_check_matrix[742] = 12'b001000110101;
    assign parity_check_matrix[743] = 12'b110111001010;
    assign parity_check_matrix[744] = 12'b010000110101;
    assign parity_check_matrix[745] = 12'b101111001010;
    assign parity_check_matrix[746] = 12'b100000110101;
    assign parity_check_matrix[747] = 12'b011111001010;
    assign parity_check_matrix[748] = 12'b000011010101;
    assign parity_check_matrix[749] = 12'b111100101010;
    assign parity_check_matrix[750] = 12'b000101010101;
    assign parity_check_matrix[751] = 12'b111010101010;
    assign parity_check_matrix[752] = 12'b001001010101;
    assign parity_check_matrix[753] = 12'b110110101010;
    assign parity_check_matrix[754] = 12'b010001010101;
    assign parity_check_matrix[755] = 12'b101110101010;
    assign parity_check_matrix[756] = 12'b100001010101;
    assign parity_check_matrix[757] = 12'b011110101010;
    assign parity_check_matrix[758] = 12'b000110010101;
    assign parity_check_matrix[759] = 12'b111001101010;
    assign parity_check_matrix[760] = 12'b001010010101;
    assign parity_check_matrix[761] = 12'b110101101010;
    assign parity_check_matrix[762] = 12'b010010010101;
    assign parity_check_matrix[763] = 12'b101101101010;
    assign parity_check_matrix[764] = 12'b100010010101;
    assign parity_check_matrix[765] = 12'b011101101010;
    assign parity_check_matrix[766] = 12'b001100010101;
    assign parity_check_matrix[767] = 12'b110011101010;
    assign parity_check_matrix[768] = 12'b010100010101;
    assign parity_check_matrix[769] = 12'b101011101010;
    assign parity_check_matrix[770] = 12'b100100010101;
    assign parity_check_matrix[771] = 12'b011011101010;
    assign parity_check_matrix[772] = 12'b011000010101;
    assign parity_check_matrix[773] = 12'b100111101010;
    assign parity_check_matrix[774] = 12'b101000010101;
    assign parity_check_matrix[775] = 12'b010111101010;
    assign parity_check_matrix[776] = 12'b110000010101;
    assign parity_check_matrix[777] = 12'b001111101010;
    assign parity_check_matrix[778] = 12'b000011100101;
    assign parity_check_matrix[779] = 12'b111100011010;
    assign parity_check_matrix[780] = 12'b000101100101;
    assign parity_check_matrix[781] = 12'b111010011010;
    assign parity_check_matrix[782] = 12'b001001100101;
    assign parity_check_matrix[783] = 12'b110110011010;
    assign parity_check_matrix[784] = 12'b010001100101;
    assign parity_check_matrix[785] = 12'b101110011010;
    assign parity_check_matrix[786] = 12'b100001100101;
    assign parity_check_matrix[787] = 12'b011110011010;
    assign parity_check_matrix[788] = 12'b000110100101;
    assign parity_check_matrix[789] = 12'b111001011010;
    assign parity_check_matrix[790] = 12'b001010100101;
    assign parity_check_matrix[791] = 12'b110101011010;
    assign parity_check_matrix[792] = 12'b010010100101;
    assign parity_check_matrix[793] = 12'b101101011010;
    assign parity_check_matrix[794] = 12'b100010100101;
    assign parity_check_matrix[795] = 12'b011101011010;
    assign parity_check_matrix[796] = 12'b001100100101;
    assign parity_check_matrix[797] = 12'b110011011010;
    assign parity_check_matrix[798] = 12'b010100100101;
    assign parity_check_matrix[799] = 12'b101011011010;
    assign parity_check_matrix[800] = 12'b100100100101;
    assign parity_check_matrix[801] = 12'b011011011010;
    assign parity_check_matrix[802] = 12'b011000100101;
    assign parity_check_matrix[803] = 12'b100111011010;
    assign parity_check_matrix[804] = 12'b101000100101;
    assign parity_check_matrix[805] = 12'b010111011010;
    assign parity_check_matrix[806] = 12'b110000100101;
    assign parity_check_matrix[807] = 12'b001111011010;
    assign parity_check_matrix[808] = 12'b000111000101;
    assign parity_check_matrix[809] = 12'b111000111010;
    assign parity_check_matrix[810] = 12'b001011000101;
    assign parity_check_matrix[811] = 12'b110100111010;
    assign parity_check_matrix[812] = 12'b010011000101;
    assign parity_check_matrix[813] = 12'b101100111010;
    assign parity_check_matrix[814] = 12'b100011000101;
    assign parity_check_matrix[815] = 12'b011100111010;
    assign parity_check_matrix[816] = 12'b001101000101;
    assign parity_check_matrix[817] = 12'b110010111010;
    assign parity_check_matrix[818] = 12'b010101000101;
    assign parity_check_matrix[819] = 12'b101010111010;
    assign parity_check_matrix[820] = 12'b100101000101;
    assign parity_check_matrix[821] = 12'b011010111010;
    assign parity_check_matrix[822] = 12'b011001000101;
    assign parity_check_matrix[823] = 12'b100110111010;
    assign parity_check_matrix[824] = 12'b101001000101;
    assign parity_check_matrix[825] = 12'b010110111010;
    assign parity_check_matrix[826] = 12'b110001000101;
    assign parity_check_matrix[827] = 12'b001110111010;
    assign parity_check_matrix[828] = 12'b001110000101;
    assign parity_check_matrix[829] = 12'b110001111010;
    assign parity_check_matrix[830] = 12'b010110000101;
    assign parity_check_matrix[831] = 12'b101001111010;
    assign parity_check_matrix[832] = 12'b100110000101;
    assign parity_check_matrix[833] = 12'b011001111010;
    assign parity_check_matrix[834] = 12'b011010000101;
    assign parity_check_matrix[835] = 12'b100101111010;
    assign parity_check_matrix[836] = 12'b101010000101;
    assign parity_check_matrix[837] = 12'b010101111010;
    assign parity_check_matrix[838] = 12'b110010000101;
    assign parity_check_matrix[839] = 12'b001101111010;
    assign parity_check_matrix[840] = 12'b011100000101;
    assign parity_check_matrix[841] = 12'b100011111010;
    assign parity_check_matrix[842] = 12'b101100000101;
    assign parity_check_matrix[843] = 12'b010011111010;
    assign parity_check_matrix[844] = 12'b110100000101;
    assign parity_check_matrix[845] = 12'b001011111010;
    assign parity_check_matrix[846] = 12'b111000000101;
    assign parity_check_matrix[847] = 12'b000111111010;
    assign parity_check_matrix[848] = 12'b000001111001;
    assign parity_check_matrix[849] = 12'b111110000110;
    assign parity_check_matrix[850] = 12'b000010111001;
    assign parity_check_matrix[851] = 12'b111101000110;
    assign parity_check_matrix[852] = 12'b000100111001;
    assign parity_check_matrix[853] = 12'b111011000110;
    assign parity_check_matrix[854] = 12'b001000111001;
    assign parity_check_matrix[855] = 12'b110111000110;
    assign parity_check_matrix[856] = 12'b010000111001;
    assign parity_check_matrix[857] = 12'b101111000110;
    assign parity_check_matrix[858] = 12'b100000111001;
    assign parity_check_matrix[859] = 12'b011111000110;
    assign parity_check_matrix[860] = 12'b000011011001;
    assign parity_check_matrix[861] = 12'b111100100110;
    assign parity_check_matrix[862] = 12'b000101011001;
    assign parity_check_matrix[863] = 12'b111010100110;
    assign parity_check_matrix[864] = 12'b001001011001;
    assign parity_check_matrix[865] = 12'b110110100110;
    assign parity_check_matrix[866] = 12'b010001011001;
    assign parity_check_matrix[867] = 12'b101110100110;
    assign parity_check_matrix[868] = 12'b100001011001;
    assign parity_check_matrix[869] = 12'b011110100110;
    assign parity_check_matrix[870] = 12'b000110011001;
    assign parity_check_matrix[871] = 12'b111001100110;
    assign parity_check_matrix[872] = 12'b001010011001;
    assign parity_check_matrix[873] = 12'b110101100110;
    assign parity_check_matrix[874] = 12'b010010011001;
    assign parity_check_matrix[875] = 12'b101101100110;
    assign parity_check_matrix[876] = 12'b100010011001;
    assign parity_check_matrix[877] = 12'b011101100110;
    assign parity_check_matrix[878] = 12'b001100011001;
    assign parity_check_matrix[879] = 12'b110011100110;
    assign parity_check_matrix[880] = 12'b010100011001;
    assign parity_check_matrix[881] = 12'b101011100110;
    assign parity_check_matrix[882] = 12'b100100011001;
    assign parity_check_matrix[883] = 12'b011011100110;
    assign parity_check_matrix[884] = 12'b011000011001;
    assign parity_check_matrix[885] = 12'b100111100110;
    assign parity_check_matrix[886] = 12'b101000011001;
    assign parity_check_matrix[887] = 12'b010111100110;
    assign parity_check_matrix[888] = 12'b110000011001;
    assign parity_check_matrix[889] = 12'b001111100110;
    assign parity_check_matrix[890] = 12'b000011101001;
    assign parity_check_matrix[891] = 12'b111100010110;
    assign parity_check_matrix[892] = 12'b000101101001;
    assign parity_check_matrix[893] = 12'b111010010110;
    assign parity_check_matrix[894] = 12'b001001101001;
    assign parity_check_matrix[895] = 12'b110110010110;
    assign parity_check_matrix[896] = 12'b010001101001;
    assign parity_check_matrix[897] = 12'b101110010110;
    assign parity_check_matrix[898] = 12'b100001101001;
    assign parity_check_matrix[899] = 12'b011110010110;
    assign parity_check_matrix[900] = 12'b000110101001;
    assign parity_check_matrix[901] = 12'b111001010110;
    assign parity_check_matrix[902] = 12'b001010101001;
    assign parity_check_matrix[903] = 12'b110101010110;
    assign parity_check_matrix[904] = 12'b010010101001;
    assign parity_check_matrix[905] = 12'b101101010110;
    assign parity_check_matrix[906] = 12'b100010101001;
    assign parity_check_matrix[907] = 12'b011101010110;
    assign parity_check_matrix[908] = 12'b001100101001;
    assign parity_check_matrix[909] = 12'b110011010110;
    assign parity_check_matrix[910] = 12'b010100101001;
    assign parity_check_matrix[911] = 12'b101011010110;
    assign parity_check_matrix[912] = 12'b100100101001;
    assign parity_check_matrix[913] = 12'b011011010110;
    assign parity_check_matrix[914] = 12'b011000101001;
    assign parity_check_matrix[915] = 12'b100111010110;
    assign parity_check_matrix[916] = 12'b101000101001;
    assign parity_check_matrix[917] = 12'b010111010110;
    assign parity_check_matrix[918] = 12'b110000101001;
    assign parity_check_matrix[919] = 12'b001111010110;
    assign parity_check_matrix[920] = 12'b000111001001;
    assign parity_check_matrix[921] = 12'b111000110110;
    assign parity_check_matrix[922] = 12'b001011001001;
    assign parity_check_matrix[923] = 12'b110100110110;
    assign parity_check_matrix[924] = 12'b010011001001;
    assign parity_check_matrix[925] = 12'b101100110110;
    assign parity_check_matrix[926] = 12'b100011001001;
    assign parity_check_matrix[927] = 12'b011100110110;
    assign parity_check_matrix[928] = 12'b001101001001;
    assign parity_check_matrix[929] = 12'b110010110110;
    assign parity_check_matrix[930] = 12'b010101001001;
    assign parity_check_matrix[931] = 12'b101010110110;
    assign parity_check_matrix[932] = 12'b100101001001;
    assign parity_check_matrix[933] = 12'b011010110110;
    assign parity_check_matrix[934] = 12'b011001001001;
    assign parity_check_matrix[935] = 12'b100110110110;
    assign parity_check_matrix[936] = 12'b101001001001;
    assign parity_check_matrix[937] = 12'b010110110110;
    assign parity_check_matrix[938] = 12'b110001001001;
    assign parity_check_matrix[939] = 12'b001110110110;
    assign parity_check_matrix[940] = 12'b001110001001;
    assign parity_check_matrix[941] = 12'b110001110110;
    assign parity_check_matrix[942] = 12'b010110001001;
    assign parity_check_matrix[943] = 12'b101001110110;
    assign parity_check_matrix[944] = 12'b100110001001;
    assign parity_check_matrix[945] = 12'b011001110110;
    assign parity_check_matrix[946] = 12'b011010001001;
    assign parity_check_matrix[947] = 12'b100101110110;
    assign parity_check_matrix[948] = 12'b101010001001;
    assign parity_check_matrix[949] = 12'b010101110110;
    assign parity_check_matrix[950] = 12'b110010001001;
    assign parity_check_matrix[951] = 12'b001101110110;
    assign parity_check_matrix[952] = 12'b011100001001;
    assign parity_check_matrix[953] = 12'b100011110110;
    assign parity_check_matrix[954] = 12'b101100001001;
    assign parity_check_matrix[955] = 12'b010011110110;
    assign parity_check_matrix[956] = 12'b110100001001;
    assign parity_check_matrix[957] = 12'b001011110110;
    assign parity_check_matrix[958] = 12'b111000001001;
    assign parity_check_matrix[959] = 12'b000111110110;
    assign parity_check_matrix[960] = 12'b000011110001;
    assign parity_check_matrix[961] = 12'b111100001110;
    assign parity_check_matrix[962] = 12'b000101110001;
    assign parity_check_matrix[963] = 12'b111010001110;
    assign parity_check_matrix[964] = 12'b001001110001;
    assign parity_check_matrix[965] = 12'b110110001110;
    assign parity_check_matrix[966] = 12'b010001110001;
    assign parity_check_matrix[967] = 12'b101110001110;
    assign parity_check_matrix[968] = 12'b100001110001;
    assign parity_check_matrix[969] = 12'b011110001110;
    assign parity_check_matrix[970] = 12'b000110110001;
    assign parity_check_matrix[971] = 12'b111001001110;
    assign parity_check_matrix[972] = 12'b001010110001;
    assign parity_check_matrix[973] = 12'b110101001110;
    assign parity_check_matrix[974] = 12'b010010110001;
    assign parity_check_matrix[975] = 12'b101101001110;
    assign parity_check_matrix[976] = 12'b100010110001;
    assign parity_check_matrix[977] = 12'b011101001110;
    assign parity_check_matrix[978] = 12'b001100110001;
    assign parity_check_matrix[979] = 12'b110011001110;
    assign parity_check_matrix[980] = 12'b010100110001;
    assign parity_check_matrix[981] = 12'b101011001110;
    assign parity_check_matrix[982] = 12'b100100110001;
    assign parity_check_matrix[983] = 12'b011011001110;
    assign parity_check_matrix[984] = 12'b011000110001;
    assign parity_check_matrix[985] = 12'b100111001110;
    assign parity_check_matrix[986] = 12'b101000110001;
    assign parity_check_matrix[987] = 12'b010111001110;
    assign parity_check_matrix[988] = 12'b110000110001;
    assign parity_check_matrix[989] = 12'b001111001110;
    assign parity_check_matrix[990] = 12'b000111010001;
    assign parity_check_matrix[991] = 12'b111000101110;
    assign parity_check_matrix[992] = 12'b001011010001;
    assign parity_check_matrix[993] = 12'b110100101110;
    assign parity_check_matrix[994] = 12'b010011010001;
    assign parity_check_matrix[995] = 12'b101100101110;
    assign parity_check_matrix[996] = 12'b100011010001;
    assign parity_check_matrix[997] = 12'b011100101110;
    assign parity_check_matrix[998] = 12'b001101010001;
    assign parity_check_matrix[999] = 12'b110010101110;
    assign parity_check_matrix[1000] = 12'b010101010001;
    assign parity_check_matrix[1001] = 12'b101010101110;
    assign parity_check_matrix[1002] = 12'b100101010001;
    assign parity_check_matrix[1003] = 12'b011010101110;
    assign parity_check_matrix[1004] = 12'b011001010001;
    assign parity_check_matrix[1005] = 12'b100110101110;
    assign parity_check_matrix[1006] = 12'b101001010001;
    assign parity_check_matrix[1007] = 12'b010110101110;
    assign parity_check_matrix[1008] = 12'b110001010001;
    assign parity_check_matrix[1009] = 12'b001110101110;
    assign parity_check_matrix[1010] = 12'b001110010001;
    assign parity_check_matrix[1011] = 12'b110001101110;
    assign parity_check_matrix[1012] = 12'b010110010001;
    assign parity_check_matrix[1013] = 12'b101001101110;
    assign parity_check_matrix[1014] = 12'b100110010001;
    assign parity_check_matrix[1015] = 12'b011001101110;
    assign parity_check_matrix[1016] = 12'b011010010001;
    assign parity_check_matrix[1017] = 12'b100101101110;
    assign parity_check_matrix[1018] = 12'b101010010001;
    assign parity_check_matrix[1019] = 12'b010101101110;
    assign parity_check_matrix[1020] = 12'b110010010001;
    assign parity_check_matrix[1021] = 12'b001101101110;
    assign parity_check_matrix[1022] = 12'b011100010001;
    assign parity_check_matrix[1023] = 12'b100011101110;
    assign parity_check_matrix[1024] = 12'b101100010001;
    assign parity_check_matrix[1025] = 12'b010011101110;
    assign parity_check_matrix[1026] = 12'b110100010001;
    assign parity_check_matrix[1027] = 12'b001011101110;
    assign parity_check_matrix[1028] = 12'b111000010001;
    assign parity_check_matrix[1029] = 12'b000111101110;
    assign parity_check_matrix[1030] = 12'b000111100001;
    assign parity_check_matrix[1031] = 12'b111000011110;
    assign parity_check_matrix[1032] = 12'b001011100001;
    assign parity_check_matrix[1033] = 12'b110100011110;
    assign parity_check_matrix[1034] = 12'b010011100001;
    assign parity_check_matrix[1035] = 12'b101100011110;
    assign parity_check_matrix[1036] = 12'b100011100001;
    assign parity_check_matrix[1037] = 12'b011100011110;
    assign parity_check_matrix[1038] = 12'b001101100001;
    assign parity_check_matrix[1039] = 12'b110010011110;
    assign parity_check_matrix[1040] = 12'b010101100001;
    assign parity_check_matrix[1041] = 12'b101010011110;
    assign parity_check_matrix[1042] = 12'b100101100001;
    assign parity_check_matrix[1043] = 12'b011010011110;
    assign parity_check_matrix[1044] = 12'b011001100001;
    assign parity_check_matrix[1045] = 12'b100110011110;
    assign parity_check_matrix[1046] = 12'b101001100001;
    assign parity_check_matrix[1047] = 12'b010110011110;
    assign parity_check_matrix[1048] = 12'b110001100001;
    assign parity_check_matrix[1049] = 12'b001110011110;
    assign parity_check_matrix[1050] = 12'b001110100001;
    assign parity_check_matrix[1051] = 12'b110001011110;
    assign parity_check_matrix[1052] = 12'b010110100001;
    assign parity_check_matrix[1053] = 12'b101001011110;
    assign parity_check_matrix[1054] = 12'b100110100001;
    assign parity_check_matrix[1055] = 12'b011001011110;
    assign parity_check_matrix[1056] = 12'b011010100001;
    assign parity_check_matrix[1057] = 12'b100101011110;
    assign parity_check_matrix[1058] = 12'b101010100001;
    assign parity_check_matrix[1059] = 12'b010101011110;
    assign parity_check_matrix[1060] = 12'b110010100001;
    assign parity_check_matrix[1061] = 12'b001101011110;
    assign parity_check_matrix[1062] = 12'b011100100001;
    assign parity_check_matrix[1063] = 12'b100011011110;
    assign parity_check_matrix[1064] = 12'b101100100001;
    assign parity_check_matrix[1065] = 12'b010011011110;
    assign parity_check_matrix[1066] = 12'b110100100001;
    assign parity_check_matrix[1067] = 12'b001011011110;
    assign parity_check_matrix[1068] = 12'b111000100001;
    assign parity_check_matrix[1069] = 12'b000111011110;
    assign parity_check_matrix[1070] = 12'b001111000001;
    assign parity_check_matrix[1071] = 12'b110000111110;
    assign parity_check_matrix[1072] = 12'b010111000001;
    assign parity_check_matrix[1073] = 12'b101000111110;
    assign parity_check_matrix[1074] = 12'b100111000001;
    assign parity_check_matrix[1075] = 12'b011000111110;
    assign parity_check_matrix[1076] = 12'b011011000001;
    assign parity_check_matrix[1077] = 12'b100100111110;
    assign parity_check_matrix[1078] = 12'b101011000001;
    assign parity_check_matrix[1079] = 12'b010100111110;
    assign parity_check_matrix[1080] = 12'b110011000001;
    assign parity_check_matrix[1081] = 12'b001100111110;
    assign parity_check_matrix[1082] = 12'b011101000001;
    assign parity_check_matrix[1083] = 12'b100010111110;
    assign parity_check_matrix[1084] = 12'b101101000001;
    assign parity_check_matrix[1085] = 12'b010010111110;
    assign parity_check_matrix[1086] = 12'b110101000001;
    assign parity_check_matrix[1087] = 12'b001010111110;
    assign parity_check_matrix[1088] = 12'b111001000001;
    assign parity_check_matrix[1089] = 12'b000110111110;
    assign parity_check_matrix[1090] = 12'b011110000001;
    assign parity_check_matrix[1091] = 12'b100001111110;
    assign parity_check_matrix[1092] = 12'b101110000001;
    assign parity_check_matrix[1093] = 12'b010001111110;
    assign parity_check_matrix[1094] = 12'b110110000001;
    assign parity_check_matrix[1095] = 12'b001001111110;
    assign parity_check_matrix[1096] = 12'b111010000001;
    assign parity_check_matrix[1097] = 12'b000101111110;
    assign parity_check_matrix[1098] = 12'b111100000001;
    assign parity_check_matrix[1099] = 12'b000011111110;
    assign parity_check_matrix[1100] = 12'b000000111110;
    assign parity_check_matrix[1101] = 12'b111111000001;
    assign parity_check_matrix[1102] = 12'b000001011110;
    assign parity_check_matrix[1103] = 12'b111110100001;
    assign parity_check_matrix[1104] = 12'b000010011110;
    assign parity_check_matrix[1105] = 12'b111101100001;
    assign parity_check_matrix[1106] = 12'b000100011110;
    assign parity_check_matrix[1107] = 12'b111011100001;
    assign parity_check_matrix[1108] = 12'b001000011110;
    assign parity_check_matrix[1109] = 12'b110111100001;
    assign parity_check_matrix[1110] = 12'b010000011110;
    assign parity_check_matrix[1111] = 12'b101111100001;
    assign parity_check_matrix[1112] = 12'b100000011110;
    assign parity_check_matrix[1113] = 12'b011111100001;
    assign parity_check_matrix[1114] = 12'b000001101110;
    assign parity_check_matrix[1115] = 12'b111110010001;
    assign parity_check_matrix[1116] = 12'b000010101110;
    assign parity_check_matrix[1117] = 12'b111101010001;
    assign parity_check_matrix[1118] = 12'b000100101110;
    assign parity_check_matrix[1119] = 12'b111011010001;
    assign parity_check_matrix[1120] = 12'b001000101110;
    assign parity_check_matrix[1121] = 12'b110111010001;
    assign parity_check_matrix[1122] = 12'b010000101110;
    assign parity_check_matrix[1123] = 12'b101111010001;
    assign parity_check_matrix[1124] = 12'b100000101110;
    assign parity_check_matrix[1125] = 12'b011111010001;
    assign parity_check_matrix[1126] = 12'b000011001110;
    assign parity_check_matrix[1127] = 12'b111100110001;
    assign parity_check_matrix[1128] = 12'b000101001110;
    assign parity_check_matrix[1129] = 12'b111010110001;
    assign parity_check_matrix[1130] = 12'b001001001110;
    assign parity_check_matrix[1131] = 12'b110110110001;
    assign parity_check_matrix[1132] = 12'b010001001110;
    assign parity_check_matrix[1133] = 12'b101110110001;
    assign parity_check_matrix[1134] = 12'b100001001110;
    assign parity_check_matrix[1135] = 12'b011110110001;
    assign parity_check_matrix[1136] = 12'b000110001110;
    assign parity_check_matrix[1137] = 12'b111001110001;
    assign parity_check_matrix[1138] = 12'b001010001110;
    assign parity_check_matrix[1139] = 12'b110101110001;
    assign parity_check_matrix[1140] = 12'b010010001110;
    assign parity_check_matrix[1141] = 12'b101101110001;
    assign parity_check_matrix[1142] = 12'b100010001110;
    assign parity_check_matrix[1143] = 12'b011101110001;
    assign parity_check_matrix[1144] = 12'b001100001110;
    assign parity_check_matrix[1145] = 12'b110011110001;
    assign parity_check_matrix[1146] = 12'b010100001110;
    assign parity_check_matrix[1147] = 12'b101011110001;
    assign parity_check_matrix[1148] = 12'b100100001110;
    assign parity_check_matrix[1149] = 12'b011011110001;
    assign parity_check_matrix[1150] = 12'b011000001110;
    assign parity_check_matrix[1151] = 12'b100111110001;
    assign parity_check_matrix[1152] = 12'b101000001110;
    assign parity_check_matrix[1153] = 12'b010111110001;
    assign parity_check_matrix[1154] = 12'b110000001110;
    assign parity_check_matrix[1155] = 12'b001111110001;
    assign parity_check_matrix[1156] = 12'b000001110110;
    assign parity_check_matrix[1157] = 12'b111110001001;
    assign parity_check_matrix[1158] = 12'b000010110110;
    assign parity_check_matrix[1159] = 12'b111101001001;
    assign parity_check_matrix[1160] = 12'b000100110110;
    assign parity_check_matrix[1161] = 12'b111011001001;
    assign parity_check_matrix[1162] = 12'b001000110110;
    assign parity_check_matrix[1163] = 12'b110111001001;
    assign parity_check_matrix[1164] = 12'b010000110110;
    assign parity_check_matrix[1165] = 12'b101111001001;
    assign parity_check_matrix[1166] = 12'b100000110110;
    assign parity_check_matrix[1167] = 12'b011111001001;
    assign parity_check_matrix[1168] = 12'b000011010110;
    assign parity_check_matrix[1169] = 12'b111100101001;
    assign parity_check_matrix[1170] = 12'b000101010110;
    assign parity_check_matrix[1171] = 12'b111010101001;
    assign parity_check_matrix[1172] = 12'b001001010110;
    assign parity_check_matrix[1173] = 12'b110110101001;
    assign parity_check_matrix[1174] = 12'b010001010110;
    assign parity_check_matrix[1175] = 12'b101110101001;
    assign parity_check_matrix[1176] = 12'b100001010110;
    assign parity_check_matrix[1177] = 12'b011110101001;
    assign parity_check_matrix[1178] = 12'b000110010110;
    assign parity_check_matrix[1179] = 12'b111001101001;
    assign parity_check_matrix[1180] = 12'b001010010110;
    assign parity_check_matrix[1181] = 12'b110101101001;
    assign parity_check_matrix[1182] = 12'b010010010110;
    assign parity_check_matrix[1183] = 12'b101101101001;
    assign parity_check_matrix[1184] = 12'b100010010110;
    assign parity_check_matrix[1185] = 12'b011101101001;
    assign parity_check_matrix[1186] = 12'b001100010110;
    assign parity_check_matrix[1187] = 12'b110011101001;
    assign parity_check_matrix[1188] = 12'b010100010110;
    assign parity_check_matrix[1189] = 12'b101011101001;
    assign parity_check_matrix[1190] = 12'b100100010110;
    assign parity_check_matrix[1191] = 12'b011011101001;
    assign parity_check_matrix[1192] = 12'b011000010110;
    assign parity_check_matrix[1193] = 12'b100111101001;
    assign parity_check_matrix[1194] = 12'b101000010110;
    assign parity_check_matrix[1195] = 12'b010111101001;
    assign parity_check_matrix[1196] = 12'b110000010110;
    assign parity_check_matrix[1197] = 12'b001111101001;
    assign parity_check_matrix[1198] = 12'b000011100110;
    assign parity_check_matrix[1199] = 12'b111100011001;
    assign parity_check_matrix[1200] = 12'b000101100110;
    assign parity_check_matrix[1201] = 12'b111010011001;
    assign parity_check_matrix[1202] = 12'b001001100110;
    assign parity_check_matrix[1203] = 12'b110110011001;
    assign parity_check_matrix[1204] = 12'b010001100110;
    assign parity_check_matrix[1205] = 12'b101110011001;
    assign parity_check_matrix[1206] = 12'b100001100110;
    assign parity_check_matrix[1207] = 12'b011110011001;
    assign parity_check_matrix[1208] = 12'b000110100110;
    assign parity_check_matrix[1209] = 12'b111001011001;
    assign parity_check_matrix[1210] = 12'b001010100110;
    assign parity_check_matrix[1211] = 12'b110101011001;
    assign parity_check_matrix[1212] = 12'b010010100110;
    assign parity_check_matrix[1213] = 12'b101101011001;
    assign parity_check_matrix[1214] = 12'b100010100110;
    assign parity_check_matrix[1215] = 12'b011101011001;
    assign parity_check_matrix[1216] = 12'b001100100110;
    assign parity_check_matrix[1217] = 12'b110011011001;
    assign parity_check_matrix[1218] = 12'b010100100110;
    assign parity_check_matrix[1219] = 12'b101011011001;
    assign parity_check_matrix[1220] = 12'b100100100110;
    assign parity_check_matrix[1221] = 12'b011011011001;
    assign parity_check_matrix[1222] = 12'b011000100110;
    assign parity_check_matrix[1223] = 12'b100111011001;
    assign parity_check_matrix[1224] = 12'b101000100110;
    assign parity_check_matrix[1225] = 12'b010111011001;
    assign parity_check_matrix[1226] = 12'b110000100110;
    assign parity_check_matrix[1227] = 12'b001111011001;
    assign parity_check_matrix[1228] = 12'b000111000110;
    assign parity_check_matrix[1229] = 12'b111000111001;
    assign parity_check_matrix[1230] = 12'b001011000110;
    assign parity_check_matrix[1231] = 12'b110100111001;
    assign parity_check_matrix[1232] = 12'b010011000110;
    assign parity_check_matrix[1233] = 12'b101100111001;
    assign parity_check_matrix[1234] = 12'b100011000110;
    assign parity_check_matrix[1235] = 12'b011100111001;
    assign parity_check_matrix[1236] = 12'b001101000110;
    assign parity_check_matrix[1237] = 12'b110010111001;
    assign parity_check_matrix[1238] = 12'b010101000110;
    assign parity_check_matrix[1239] = 12'b101010111001;
    assign parity_check_matrix[1240] = 12'b100101000110;
    assign parity_check_matrix[1241] = 12'b011010111001;
    assign parity_check_matrix[1242] = 12'b011001000110;
    assign parity_check_matrix[1243] = 12'b100110111001;
    assign parity_check_matrix[1244] = 12'b101001000110;
    assign parity_check_matrix[1245] = 12'b010110111001;
    assign parity_check_matrix[1246] = 12'b110001000110;
    assign parity_check_matrix[1247] = 12'b001110111001;
    assign parity_check_matrix[1248] = 12'b001110000110;
    assign parity_check_matrix[1249] = 12'b110001111001;
    assign parity_check_matrix[1250] = 12'b010110000110;
    assign parity_check_matrix[1251] = 12'b101001111001;
    assign parity_check_matrix[1252] = 12'b100110000110;
    assign parity_check_matrix[1253] = 12'b011001111001;
    assign parity_check_matrix[1254] = 12'b011010000110;
    assign parity_check_matrix[1255] = 12'b100101111001;
    assign parity_check_matrix[1256] = 12'b101010000110;
    assign parity_check_matrix[1257] = 12'b010101111001;
    assign parity_check_matrix[1258] = 12'b110010000110;
    assign parity_check_matrix[1259] = 12'b001101111001;
    assign parity_check_matrix[1260] = 12'b011100000110;
    assign parity_check_matrix[1261] = 12'b100011111001;
    assign parity_check_matrix[1262] = 12'b101100000110;
    assign parity_check_matrix[1263] = 12'b010011111001;
    assign parity_check_matrix[1264] = 12'b110100000110;
    assign parity_check_matrix[1265] = 12'b001011111001;
    assign parity_check_matrix[1266] = 12'b111000000110;
    assign parity_check_matrix[1267] = 12'b000111111001;
    assign parity_check_matrix[1268] = 12'b000001111010;
    assign parity_check_matrix[1269] = 12'b111110000101;
    assign parity_check_matrix[1270] = 12'b000010111010;
    assign parity_check_matrix[1271] = 12'b111101000101;
    assign parity_check_matrix[1272] = 12'b000100111010;
    assign parity_check_matrix[1273] = 12'b111011000101;
    assign parity_check_matrix[1274] = 12'b001000111010;
    assign parity_check_matrix[1275] = 12'b110111000101;
    assign parity_check_matrix[1276] = 12'b010000111010;
    assign parity_check_matrix[1277] = 12'b101111000101;
    assign parity_check_matrix[1278] = 12'b100000111010;
    assign parity_check_matrix[1279] = 12'b011111000101;
    assign parity_check_matrix[1280] = 12'b000011011010;
    assign parity_check_matrix[1281] = 12'b111100100101;
    assign parity_check_matrix[1282] = 12'b000101011010;
    assign parity_check_matrix[1283] = 12'b111010100101;
    assign parity_check_matrix[1284] = 12'b001001011010;
    assign parity_check_matrix[1285] = 12'b110110100101;
    assign parity_check_matrix[1286] = 12'b010001011010;
    assign parity_check_matrix[1287] = 12'b101110100101;
    assign parity_check_matrix[1288] = 12'b100001011010;
    assign parity_check_matrix[1289] = 12'b011110100101;
    assign parity_check_matrix[1290] = 12'b000110011010;
    assign parity_check_matrix[1291] = 12'b111001100101;
    assign parity_check_matrix[1292] = 12'b001010011010;
    assign parity_check_matrix[1293] = 12'b110101100101;
    assign parity_check_matrix[1294] = 12'b010010011010;
    assign parity_check_matrix[1295] = 12'b101101100101;
    assign parity_check_matrix[1296] = 12'b100010011010;
    assign parity_check_matrix[1297] = 12'b011101100101;
    assign parity_check_matrix[1298] = 12'b001100011010;
    assign parity_check_matrix[1299] = 12'b110011100101;
    assign parity_check_matrix[1300] = 12'b010100011010;
    assign parity_check_matrix[1301] = 12'b101011100101;
    assign parity_check_matrix[1302] = 12'b100100011010;
    assign parity_check_matrix[1303] = 12'b011011100101;
    assign parity_check_matrix[1304] = 12'b011000011010;
    assign parity_check_matrix[1305] = 12'b100111100101;
    assign parity_check_matrix[1306] = 12'b101000011010;
    assign parity_check_matrix[1307] = 12'b010111100101;
    assign parity_check_matrix[1308] = 12'b110000011010;
    assign parity_check_matrix[1309] = 12'b001111100101;
    assign parity_check_matrix[1310] = 12'b000011101010;
    assign parity_check_matrix[1311] = 12'b111100010101;
    assign parity_check_matrix[1312] = 12'b000101101010;
    assign parity_check_matrix[1313] = 12'b111010010101;
    assign parity_check_matrix[1314] = 12'b001001101010;
    assign parity_check_matrix[1315] = 12'b110110010101;
    assign parity_check_matrix[1316] = 12'b010001101010;
    assign parity_check_matrix[1317] = 12'b101110010101;
    assign parity_check_matrix[1318] = 12'b100001101010;
    assign parity_check_matrix[1319] = 12'b011110010101;
    assign parity_check_matrix[1320] = 12'b000110101010;
    assign parity_check_matrix[1321] = 12'b111001010101;
    assign parity_check_matrix[1322] = 12'b001010101010;
    assign parity_check_matrix[1323] = 12'b110101010101;
    assign parity_check_matrix[1324] = 12'b010010101010;
    assign parity_check_matrix[1325] = 12'b101101010101;
    assign parity_check_matrix[1326] = 12'b100010101010;
    assign parity_check_matrix[1327] = 12'b011101010101;
    assign parity_check_matrix[1328] = 12'b001100101010;
    assign parity_check_matrix[1329] = 12'b110011010101;
    assign parity_check_matrix[1330] = 12'b010100101010;
    assign parity_check_matrix[1331] = 12'b101011010101;
    assign parity_check_matrix[1332] = 12'b100100101010;
    assign parity_check_matrix[1333] = 12'b011011010101;
    assign parity_check_matrix[1334] = 12'b011000101010;
    assign parity_check_matrix[1335] = 12'b100111010101;
    assign parity_check_matrix[1336] = 12'b101000101010;
    assign parity_check_matrix[1337] = 12'b010111010101;
    assign parity_check_matrix[1338] = 12'b110000101010;
    assign parity_check_matrix[1339] = 12'b001111010101;
    assign parity_check_matrix[1340] = 12'b000111001010;
    assign parity_check_matrix[1341] = 12'b111000110101;
    assign parity_check_matrix[1342] = 12'b001011001010;
    assign parity_check_matrix[1343] = 12'b110100110101;
    assign parity_check_matrix[1344] = 12'b010011001010;
    assign parity_check_matrix[1345] = 12'b101100110101;
    assign parity_check_matrix[1346] = 12'b100011001010;
    assign parity_check_matrix[1347] = 12'b011100110101;
    assign parity_check_matrix[1348] = 12'b001101001010;
    assign parity_check_matrix[1349] = 12'b110010110101;
    assign parity_check_matrix[1350] = 12'b010101001010;
    assign parity_check_matrix[1351] = 12'b101010110101;
    assign parity_check_matrix[1352] = 12'b100101001010;
    assign parity_check_matrix[1353] = 12'b011010110101;
    assign parity_check_matrix[1354] = 12'b011001001010;
    assign parity_check_matrix[1355] = 12'b100110110101;
    assign parity_check_matrix[1356] = 12'b101001001010;
    assign parity_check_matrix[1357] = 12'b010110110101;
    assign parity_check_matrix[1358] = 12'b110001001010;
    assign parity_check_matrix[1359] = 12'b001110110101;
    assign parity_check_matrix[1360] = 12'b001110001010;
    assign parity_check_matrix[1361] = 12'b110001110101;
    assign parity_check_matrix[1362] = 12'b010110001010;
    assign parity_check_matrix[1363] = 12'b101001110101;
    assign parity_check_matrix[1364] = 12'b100110001010;
    assign parity_check_matrix[1365] = 12'b011001110101;
    assign parity_check_matrix[1366] = 12'b011010001010;
    assign parity_check_matrix[1367] = 12'b100101110101;
    assign parity_check_matrix[1368] = 12'b101010001010;
    assign parity_check_matrix[1369] = 12'b010101110101;
    assign parity_check_matrix[1370] = 12'b110010001010;
    assign parity_check_matrix[1371] = 12'b001101110101;
    assign parity_check_matrix[1372] = 12'b011100001010;
    assign parity_check_matrix[1373] = 12'b100011110101;
    assign parity_check_matrix[1374] = 12'b101100001010;
    assign parity_check_matrix[1375] = 12'b010011110101;
    assign parity_check_matrix[1376] = 12'b110100001010;
    assign parity_check_matrix[1377] = 12'b001011110101;
    assign parity_check_matrix[1378] = 12'b111000001010;
    assign parity_check_matrix[1379] = 12'b000111110101;
    assign parity_check_matrix[1380] = 12'b000011110010;
    assign parity_check_matrix[1381] = 12'b111100001101;
    assign parity_check_matrix[1382] = 12'b000101110010;
    assign parity_check_matrix[1383] = 12'b111010001101;
    assign parity_check_matrix[1384] = 12'b001001110010;
    assign parity_check_matrix[1385] = 12'b110110001101;
    assign parity_check_matrix[1386] = 12'b010001110010;
    assign parity_check_matrix[1387] = 12'b101110001101;
    assign parity_check_matrix[1388] = 12'b100001110010;
    assign parity_check_matrix[1389] = 12'b011110001101;
    assign parity_check_matrix[1390] = 12'b000110110010;
    assign parity_check_matrix[1391] = 12'b111001001101;
    assign parity_check_matrix[1392] = 12'b001010110010;
    assign parity_check_matrix[1393] = 12'b110101001101;
    assign parity_check_matrix[1394] = 12'b010010110010;
    assign parity_check_matrix[1395] = 12'b101101001101;
    assign parity_check_matrix[1396] = 12'b100010110010;
    assign parity_check_matrix[1397] = 12'b011101001101;
    assign parity_check_matrix[1398] = 12'b001100110010;
    assign parity_check_matrix[1399] = 12'b110011001101;
    assign parity_check_matrix[1400] = 12'b010100110010;
    assign parity_check_matrix[1401] = 12'b101011001101;
    assign parity_check_matrix[1402] = 12'b100100110010;
    assign parity_check_matrix[1403] = 12'b011011001101;
    assign parity_check_matrix[1404] = 12'b011000110010;
    assign parity_check_matrix[1405] = 12'b100111001101;
    assign parity_check_matrix[1406] = 12'b101000110010;
    assign parity_check_matrix[1407] = 12'b010111001101;
    assign parity_check_matrix[1408] = 12'b110000110010;
    assign parity_check_matrix[1409] = 12'b001111001101;
    assign parity_check_matrix[1410] = 12'b000111010010;
    assign parity_check_matrix[1411] = 12'b111000101101;
    assign parity_check_matrix[1412] = 12'b001011010010;
    assign parity_check_matrix[1413] = 12'b110100101101;
    assign parity_check_matrix[1414] = 12'b010011010010;
    assign parity_check_matrix[1415] = 12'b101100101101;
    assign parity_check_matrix[1416] = 12'b100011010010;
    assign parity_check_matrix[1417] = 12'b011100101101;
    assign parity_check_matrix[1418] = 12'b001101010010;
    assign parity_check_matrix[1419] = 12'b110010101101;
    assign parity_check_matrix[1420] = 12'b010101010010;
    assign parity_check_matrix[1421] = 12'b101010101101;
    assign parity_check_matrix[1422] = 12'b100101010010;
    assign parity_check_matrix[1423] = 12'b011010101101;
    assign parity_check_matrix[1424] = 12'b011001010010;
    assign parity_check_matrix[1425] = 12'b100110101101;
    assign parity_check_matrix[1426] = 12'b101001010010;
    assign parity_check_matrix[1427] = 12'b010110101101;
    assign parity_check_matrix[1428] = 12'b110001010010;
    assign parity_check_matrix[1429] = 12'b001110101101;
    assign parity_check_matrix[1430] = 12'b001110010010;
    assign parity_check_matrix[1431] = 12'b110001101101;
    assign parity_check_matrix[1432] = 12'b010110010010;
    assign parity_check_matrix[1433] = 12'b101001101101;
    assign parity_check_matrix[1434] = 12'b100110010010;
    assign parity_check_matrix[1435] = 12'b011001101101;
    assign parity_check_matrix[1436] = 12'b011010010010;
    assign parity_check_matrix[1437] = 12'b100101101101;
    assign parity_check_matrix[1438] = 12'b101010010010;
    assign parity_check_matrix[1439] = 12'b010101101101;
    assign parity_check_matrix[1440] = 12'b110010010010;
    assign parity_check_matrix[1441] = 12'b001101101101;
    assign parity_check_matrix[1442] = 12'b011100010010;
    assign parity_check_matrix[1443] = 12'b100011101101;
    assign parity_check_matrix[1444] = 12'b101100010010;
    assign parity_check_matrix[1445] = 12'b010011101101;
    assign parity_check_matrix[1446] = 12'b110100010010;
    assign parity_check_matrix[1447] = 12'b001011101101;
    assign parity_check_matrix[1448] = 12'b111000010010;
    assign parity_check_matrix[1449] = 12'b000111101101;
    assign parity_check_matrix[1450] = 12'b000111100010;
    assign parity_check_matrix[1451] = 12'b111000011101;
    assign parity_check_matrix[1452] = 12'b001011100010;
    assign parity_check_matrix[1453] = 12'b110100011101;
    assign parity_check_matrix[1454] = 12'b010011100010;
    assign parity_check_matrix[1455] = 12'b101100011101;
    assign parity_check_matrix[1456] = 12'b100011100010;
    assign parity_check_matrix[1457] = 12'b011100011101;
    assign parity_check_matrix[1458] = 12'b001101100010;
    assign parity_check_matrix[1459] = 12'b110010011101;
    assign parity_check_matrix[1460] = 12'b010101100010;
    assign parity_check_matrix[1461] = 12'b101010011101;
    assign parity_check_matrix[1462] = 12'b100101100010;
    assign parity_check_matrix[1463] = 12'b011010011101;
    assign parity_check_matrix[1464] = 12'b011001100010;
    assign parity_check_matrix[1465] = 12'b100110011101;
    assign parity_check_matrix[1466] = 12'b101001100010;
    assign parity_check_matrix[1467] = 12'b010110011101;
    assign parity_check_matrix[1468] = 12'b110001100010;
    assign parity_check_matrix[1469] = 12'b001110011101;
    assign parity_check_matrix[1470] = 12'b001110100010;
    assign parity_check_matrix[1471] = 12'b110001011101;
    assign parity_check_matrix[1472] = 12'b010110100010;
    assign parity_check_matrix[1473] = 12'b101001011101;
    assign parity_check_matrix[1474] = 12'b100110100010;
    assign parity_check_matrix[1475] = 12'b011001011101;
    assign parity_check_matrix[1476] = 12'b011010100010;
    assign parity_check_matrix[1477] = 12'b100101011101;
    assign parity_check_matrix[1478] = 12'b101010100010;
    assign parity_check_matrix[1479] = 12'b010101011101;
    assign parity_check_matrix[1480] = 12'b110010100010;
    assign parity_check_matrix[1481] = 12'b001101011101;
    assign parity_check_matrix[1482] = 12'b011100100010;
    assign parity_check_matrix[1483] = 12'b100011011101;
    assign parity_check_matrix[1484] = 12'b101100100010;
    assign parity_check_matrix[1485] = 12'b010011011101;
    assign parity_check_matrix[1486] = 12'b110100100010;
    assign parity_check_matrix[1487] = 12'b001011011101;
    assign parity_check_matrix[1488] = 12'b111000100010;
    assign parity_check_matrix[1489] = 12'b000111011101;
    assign parity_check_matrix[1490] = 12'b001111000010;
    assign parity_check_matrix[1491] = 12'b110000111101;
    assign parity_check_matrix[1492] = 12'b010111000010;
    assign parity_check_matrix[1493] = 12'b101000111101;
    assign parity_check_matrix[1494] = 12'b100111000010;
    assign parity_check_matrix[1495] = 12'b011000111101;
    assign parity_check_matrix[1496] = 12'b011011000010;
    assign parity_check_matrix[1497] = 12'b100100111101;
    assign parity_check_matrix[1498] = 12'b101011000010;
    assign parity_check_matrix[1499] = 12'b010100111101;
    assign parity_check_matrix[1500] = 12'b110011000010;
    assign parity_check_matrix[1501] = 12'b001100111101;
    assign parity_check_matrix[1502] = 12'b011101000010;
    assign parity_check_matrix[1503] = 12'b100010111101;
    assign parity_check_matrix[1504] = 12'b101101000010;
    assign parity_check_matrix[1505] = 12'b010010111101;
    assign parity_check_matrix[1506] = 12'b110101000010;
    assign parity_check_matrix[1507] = 12'b001010111101;
    assign parity_check_matrix[1508] = 12'b111001000010;
    assign parity_check_matrix[1509] = 12'b000110111101;
    assign parity_check_matrix[1510] = 12'b011110000010;
    assign parity_check_matrix[1511] = 12'b100001111101;
    assign parity_check_matrix[1512] = 12'b101110000010;
    assign parity_check_matrix[1513] = 12'b010001111101;
    assign parity_check_matrix[1514] = 12'b110110000010;
    assign parity_check_matrix[1515] = 12'b001001111101;
    assign parity_check_matrix[1516] = 12'b111010000010;
    assign parity_check_matrix[1517] = 12'b000101111101;
    assign parity_check_matrix[1518] = 12'b111100000010;
    assign parity_check_matrix[1519] = 12'b000011111101;
    assign parity_check_matrix[1520] = 12'b000001111100;
    assign parity_check_matrix[1521] = 12'b111110000011;
    assign parity_check_matrix[1522] = 12'b000010111100;
    assign parity_check_matrix[1523] = 12'b111101000011;
    assign parity_check_matrix[1524] = 12'b000100111100;
    assign parity_check_matrix[1525] = 12'b111011000011;
    assign parity_check_matrix[1526] = 12'b001000111100;
    assign parity_check_matrix[1527] = 12'b110111000011;
    assign parity_check_matrix[1528] = 12'b010000111100;
    assign parity_check_matrix[1529] = 12'b101111000011;
    assign parity_check_matrix[1530] = 12'b100000111100;
    assign parity_check_matrix[1531] = 12'b011111000011;
    assign parity_check_matrix[1532] = 12'b000011011100;
    assign parity_check_matrix[1533] = 12'b111100100011;
    assign parity_check_matrix[1534] = 12'b000101011100;
    assign parity_check_matrix[1535] = 12'b111010100011;
    assign parity_check_matrix[1536] = 12'b001001011100;
    assign parity_check_matrix[1537] = 12'b110110100011;
    assign parity_check_matrix[1538] = 12'b010001011100;
    assign parity_check_matrix[1539] = 12'b101110100011;
    assign parity_check_matrix[1540] = 12'b100001011100;
    assign parity_check_matrix[1541] = 12'b011110100011;
    assign parity_check_matrix[1542] = 12'b000110011100;
    assign parity_check_matrix[1543] = 12'b111001100011;
    assign parity_check_matrix[1544] = 12'b001010011100;
    assign parity_check_matrix[1545] = 12'b110101100011;
    assign parity_check_matrix[1546] = 12'b010010011100;
    assign parity_check_matrix[1547] = 12'b101101100011;
    assign parity_check_matrix[1548] = 12'b100010011100;
    assign parity_check_matrix[1549] = 12'b011101100011;
    assign parity_check_matrix[1550] = 12'b001100011100;
    assign parity_check_matrix[1551] = 12'b110011100011;
    assign parity_check_matrix[1552] = 12'b010100011100;
    assign parity_check_matrix[1553] = 12'b101011100011;
    assign parity_check_matrix[1554] = 12'b100100011100;
    assign parity_check_matrix[1555] = 12'b011011100011;
    assign parity_check_matrix[1556] = 12'b011000011100;
    assign parity_check_matrix[1557] = 12'b100111100011;
    assign parity_check_matrix[1558] = 12'b101000011100;
    assign parity_check_matrix[1559] = 12'b010111100011;
    assign parity_check_matrix[1560] = 12'b110000011100;
    assign parity_check_matrix[1561] = 12'b001111100011;
    assign parity_check_matrix[1562] = 12'b000011101100;
    assign parity_check_matrix[1563] = 12'b111100010011;
    assign parity_check_matrix[1564] = 12'b000101101100;
    assign parity_check_matrix[1565] = 12'b111010010011;
    assign parity_check_matrix[1566] = 12'b001001101100;
    assign parity_check_matrix[1567] = 12'b110110010011;
    assign parity_check_matrix[1568] = 12'b010001101100;
    assign parity_check_matrix[1569] = 12'b101110010011;
    assign parity_check_matrix[1570] = 12'b100001101100;
    assign parity_check_matrix[1571] = 12'b011110010011;
    assign parity_check_matrix[1572] = 12'b000110101100;
    assign parity_check_matrix[1573] = 12'b111001010011;
    assign parity_check_matrix[1574] = 12'b001010101100;
    assign parity_check_matrix[1575] = 12'b110101010011;
    assign parity_check_matrix[1576] = 12'b010010101100;
    assign parity_check_matrix[1577] = 12'b101101010011;
    assign parity_check_matrix[1578] = 12'b100010101100;
    assign parity_check_matrix[1579] = 12'b011101010011;
    assign parity_check_matrix[1580] = 12'b001100101100;
    assign parity_check_matrix[1581] = 12'b110011010011;
    assign parity_check_matrix[1582] = 12'b010100101100;
    assign parity_check_matrix[1583] = 12'b101011010011;
    assign parity_check_matrix[1584] = 12'b100100101100;
    assign parity_check_matrix[1585] = 12'b011011010011;
    assign parity_check_matrix[1586] = 12'b011000101100;
    assign parity_check_matrix[1587] = 12'b100111010011;
    assign parity_check_matrix[1588] = 12'b101000101100;
    assign parity_check_matrix[1589] = 12'b010111010011;
    assign parity_check_matrix[1590] = 12'b110000101100;
    assign parity_check_matrix[1591] = 12'b001111010011;
    assign parity_check_matrix[1592] = 12'b000111001100;
    assign parity_check_matrix[1593] = 12'b111000110011;
    assign parity_check_matrix[1594] = 12'b001011001100;
    assign parity_check_matrix[1595] = 12'b110100110011;
    assign parity_check_matrix[1596] = 12'b010011001100;
    assign parity_check_matrix[1597] = 12'b101100110011;
    assign parity_check_matrix[1598] = 12'b100011001100;
    assign parity_check_matrix[1599] = 12'b011100110011;
    assign parity_check_matrix[1600] = 12'b001101001100;
    assign parity_check_matrix[1601] = 12'b110010110011;
    assign parity_check_matrix[1602] = 12'b010101001100;
    assign parity_check_matrix[1603] = 12'b101010110011;
    assign parity_check_matrix[1604] = 12'b100101001100;
    assign parity_check_matrix[1605] = 12'b011010110011;
    assign parity_check_matrix[1606] = 12'b011001001100;
    assign parity_check_matrix[1607] = 12'b100110110011;
    assign parity_check_matrix[1608] = 12'b101001001100;
    assign parity_check_matrix[1609] = 12'b010110110011;
    assign parity_check_matrix[1610] = 12'b110001001100;
    assign parity_check_matrix[1611] = 12'b001110110011;
    assign parity_check_matrix[1612] = 12'b001110001100;
    assign parity_check_matrix[1613] = 12'b110001110011;
    assign parity_check_matrix[1614] = 12'b010110001100;
    assign parity_check_matrix[1615] = 12'b101001110011;
    assign parity_check_matrix[1616] = 12'b100110001100;
    assign parity_check_matrix[1617] = 12'b011001110011;
    assign parity_check_matrix[1618] = 12'b011010001100;
    assign parity_check_matrix[1619] = 12'b100101110011;
    assign parity_check_matrix[1620] = 12'b101010001100;
    assign parity_check_matrix[1621] = 12'b010101110011;
    assign parity_check_matrix[1622] = 12'b110010001100;
    assign parity_check_matrix[1623] = 12'b001101110011;
    assign parity_check_matrix[1624] = 12'b011100001100;
    assign parity_check_matrix[1625] = 12'b100011110011;
    assign parity_check_matrix[1626] = 12'b101100001100;
    assign parity_check_matrix[1627] = 12'b010011110011;
    assign parity_check_matrix[1628] = 12'b110100001100;
    assign parity_check_matrix[1629] = 12'b001011110011;
    assign parity_check_matrix[1630] = 12'b111000001100;
    assign parity_check_matrix[1631] = 12'b000111110011;
    assign parity_check_matrix[1632] = 12'b000011110100;
    assign parity_check_matrix[1633] = 12'b111100001011;
    assign parity_check_matrix[1634] = 12'b000101110100;
    assign parity_check_matrix[1635] = 12'b111010001011;
    assign parity_check_matrix[1636] = 12'b001001110100;
    assign parity_check_matrix[1637] = 12'b110110001011;
    assign parity_check_matrix[1638] = 12'b010001110100;
    assign parity_check_matrix[1639] = 12'b101110001011;
    assign parity_check_matrix[1640] = 12'b100001110100;
    assign parity_check_matrix[1641] = 12'b011110001011;
    assign parity_check_matrix[1642] = 12'b000110110100;
    assign parity_check_matrix[1643] = 12'b111001001011;
    assign parity_check_matrix[1644] = 12'b001010110100;
    assign parity_check_matrix[1645] = 12'b110101001011;
    assign parity_check_matrix[1646] = 12'b010010110100;
    assign parity_check_matrix[1647] = 12'b101101001011;
    assign parity_check_matrix[1648] = 12'b100010110100;
    assign parity_check_matrix[1649] = 12'b011101001011;
    assign parity_check_matrix[1650] = 12'b001100110100;
    assign parity_check_matrix[1651] = 12'b110011001011;
    assign parity_check_matrix[1652] = 12'b010100110100;
    assign parity_check_matrix[1653] = 12'b101011001011;
    assign parity_check_matrix[1654] = 12'b100100110100;
    assign parity_check_matrix[1655] = 12'b011011001011;
    assign parity_check_matrix[1656] = 12'b011000110100;
    assign parity_check_matrix[1657] = 12'b100111001011;
    assign parity_check_matrix[1658] = 12'b101000110100;
    assign parity_check_matrix[1659] = 12'b010111001011;
    assign parity_check_matrix[1660] = 12'b110000110100;
    assign parity_check_matrix[1661] = 12'b001111001011;
    assign parity_check_matrix[1662] = 12'b000111010100;
    assign parity_check_matrix[1663] = 12'b111000101011;
    assign parity_check_matrix[1664] = 12'b001011010100;
    assign parity_check_matrix[1665] = 12'b110100101011;
    assign parity_check_matrix[1666] = 12'b010011010100;
    assign parity_check_matrix[1667] = 12'b101100101011;
    assign parity_check_matrix[1668] = 12'b100011010100;
    assign parity_check_matrix[1669] = 12'b011100101011;
    assign parity_check_matrix[1670] = 12'b001101010100;
    assign parity_check_matrix[1671] = 12'b110010101011;
    assign parity_check_matrix[1672] = 12'b010101010100;
    assign parity_check_matrix[1673] = 12'b101010101011;
    assign parity_check_matrix[1674] = 12'b100101010100;
    assign parity_check_matrix[1675] = 12'b011010101011;
    assign parity_check_matrix[1676] = 12'b011001010100;
    assign parity_check_matrix[1677] = 12'b100110101011;
    assign parity_check_matrix[1678] = 12'b101001010100;
    assign parity_check_matrix[1679] = 12'b010110101011;
    assign parity_check_matrix[1680] = 12'b110001010100;
    assign parity_check_matrix[1681] = 12'b001110101011;
    assign parity_check_matrix[1682] = 12'b001110010100;
    assign parity_check_matrix[1683] = 12'b110001101011;
    assign parity_check_matrix[1684] = 12'b010110010100;
    assign parity_check_matrix[1685] = 12'b101001101011;
    assign parity_check_matrix[1686] = 12'b100110010100;
    assign parity_check_matrix[1687] = 12'b011001101011;
    assign parity_check_matrix[1688] = 12'b011010010100;
    assign parity_check_matrix[1689] = 12'b100101101011;
    assign parity_check_matrix[1690] = 12'b101010010100;
    assign parity_check_matrix[1691] = 12'b010101101011;
    assign parity_check_matrix[1692] = 12'b110010010100;
    assign parity_check_matrix[1693] = 12'b001101101011;
    assign parity_check_matrix[1694] = 12'b011100010100;
    assign parity_check_matrix[1695] = 12'b100011101011;
    assign parity_check_matrix[1696] = 12'b101100010100;
    assign parity_check_matrix[1697] = 12'b010011101011;
    assign parity_check_matrix[1698] = 12'b110100010100;
    assign parity_check_matrix[1699] = 12'b001011101011;
    assign parity_check_matrix[1700] = 12'b111000010100;
    assign parity_check_matrix[1701] = 12'b000111101011;
    assign parity_check_matrix[1702] = 12'b000111100100;
    assign parity_check_matrix[1703] = 12'b111000011011;
    assign parity_check_matrix[1704] = 12'b001011100100;
    assign parity_check_matrix[1705] = 12'b110100011011;
    assign parity_check_matrix[1706] = 12'b010011100100;
    assign parity_check_matrix[1707] = 12'b101100011011;
    assign parity_check_matrix[1708] = 12'b100011100100;
    assign parity_check_matrix[1709] = 12'b011100011011;
    assign parity_check_matrix[1710] = 12'b001101100100;
    assign parity_check_matrix[1711] = 12'b110010011011;
    assign parity_check_matrix[1712] = 12'b010101100100;
    assign parity_check_matrix[1713] = 12'b101010011011;
    assign parity_check_matrix[1714] = 12'b100101100100;
    assign parity_check_matrix[1715] = 12'b011010011011;
    assign parity_check_matrix[1716] = 12'b011001100100;
    assign parity_check_matrix[1717] = 12'b100110011011;
    assign parity_check_matrix[1718] = 12'b101001100100;
    assign parity_check_matrix[1719] = 12'b010110011011;
    assign parity_check_matrix[1720] = 12'b110001100100;
    assign parity_check_matrix[1721] = 12'b001110011011;
    assign parity_check_matrix[1722] = 12'b001110100100;
    assign parity_check_matrix[1723] = 12'b110001011011;
    assign parity_check_matrix[1724] = 12'b010110100100;
    assign parity_check_matrix[1725] = 12'b101001011011;
    assign parity_check_matrix[1726] = 12'b100110100100;
    assign parity_check_matrix[1727] = 12'b011001011011;
    assign parity_check_matrix[1728] = 12'b011010100100;
    assign parity_check_matrix[1729] = 12'b100101011011;
    assign parity_check_matrix[1730] = 12'b101010100100;
    assign parity_check_matrix[1731] = 12'b010101011011;
    assign parity_check_matrix[1732] = 12'b110010100100;
    assign parity_check_matrix[1733] = 12'b001101011011;
    assign parity_check_matrix[1734] = 12'b011100100100;
    assign parity_check_matrix[1735] = 12'b100011011011;
    assign parity_check_matrix[1736] = 12'b101100100100;
    assign parity_check_matrix[1737] = 12'b010011011011;
    assign parity_check_matrix[1738] = 12'b110100100100;
    assign parity_check_matrix[1739] = 12'b001011011011;
    assign parity_check_matrix[1740] = 12'b111000100100;
    assign parity_check_matrix[1741] = 12'b000111011011;
    assign parity_check_matrix[1742] = 12'b001111000100;
    assign parity_check_matrix[1743] = 12'b110000111011;
    assign parity_check_matrix[1744] = 12'b010111000100;
    assign parity_check_matrix[1745] = 12'b101000111011;
    assign parity_check_matrix[1746] = 12'b100111000100;
    assign parity_check_matrix[1747] = 12'b011000111011;
    assign parity_check_matrix[1748] = 12'b011011000100;
    assign parity_check_matrix[1749] = 12'b100100111011;
    assign parity_check_matrix[1750] = 12'b101011000100;
    assign parity_check_matrix[1751] = 12'b010100111011;
    assign parity_check_matrix[1752] = 12'b110011000100;
    assign parity_check_matrix[1753] = 12'b001100111011;
    assign parity_check_matrix[1754] = 12'b011101000100;
    assign parity_check_matrix[1755] = 12'b100010111011;
    assign parity_check_matrix[1756] = 12'b101101000100;
    assign parity_check_matrix[1757] = 12'b010010111011;
    assign parity_check_matrix[1758] = 12'b110101000100;
    assign parity_check_matrix[1759] = 12'b001010111011;
    assign parity_check_matrix[1760] = 12'b111001000100;
    assign parity_check_matrix[1761] = 12'b000110111011;
    assign parity_check_matrix[1762] = 12'b011110000100;
    assign parity_check_matrix[1763] = 12'b100001111011;
    assign parity_check_matrix[1764] = 12'b101110000100;
    assign parity_check_matrix[1765] = 12'b010001111011;
    assign parity_check_matrix[1766] = 12'b110110000100;
    assign parity_check_matrix[1767] = 12'b001001111011;
    assign parity_check_matrix[1768] = 12'b111010000100;
    assign parity_check_matrix[1769] = 12'b000101111011;
    assign parity_check_matrix[1770] = 12'b111100000100;
    assign parity_check_matrix[1771] = 12'b000011111011;
    assign parity_check_matrix[1772] = 12'b000011111000;
    assign parity_check_matrix[1773] = 12'b111100000111;
    assign parity_check_matrix[1774] = 12'b000101111000;
    assign parity_check_matrix[1775] = 12'b111010000111;
    assign parity_check_matrix[1776] = 12'b001001111000;
    assign parity_check_matrix[1777] = 12'b110110000111;
    assign parity_check_matrix[1778] = 12'b010001111000;
    assign parity_check_matrix[1779] = 12'b101110000111;
    assign parity_check_matrix[1780] = 12'b100001111000;
    assign parity_check_matrix[1781] = 12'b011110000111;
    assign parity_check_matrix[1782] = 12'b000110111000;
    assign parity_check_matrix[1783] = 12'b111001000111;
    assign parity_check_matrix[1784] = 12'b001010111000;
    assign parity_check_matrix[1785] = 12'b110101000111;
    assign parity_check_matrix[1786] = 12'b010010111000;
    assign parity_check_matrix[1787] = 12'b101101000111;
    assign parity_check_matrix[1788] = 12'b100010111000;
    assign parity_check_matrix[1789] = 12'b011101000111;
    assign parity_check_matrix[1790] = 12'b001100111000;
    assign parity_check_matrix[1791] = 12'b110011000111;
    assign parity_check_matrix[1792] = 12'b010100111000;
    assign parity_check_matrix[1793] = 12'b101011000111;
    assign parity_check_matrix[1794] = 12'b100100111000;
    assign parity_check_matrix[1795] = 12'b011011000111;
    assign parity_check_matrix[1796] = 12'b011000111000;
    assign parity_check_matrix[1797] = 12'b100111000111;
    assign parity_check_matrix[1798] = 12'b101000111000;
    assign parity_check_matrix[1799] = 12'b010111000111;
    assign parity_check_matrix[1800] = 12'b110000111000;
    assign parity_check_matrix[1801] = 12'b001111000111;
    assign parity_check_matrix[1802] = 12'b000111011000;
    assign parity_check_matrix[1803] = 12'b111000100111;
    assign parity_check_matrix[1804] = 12'b001011011000;
    assign parity_check_matrix[1805] = 12'b110100100111;
    assign parity_check_matrix[1806] = 12'b010011011000;
    assign parity_check_matrix[1807] = 12'b101100100111;
    assign parity_check_matrix[1808] = 12'b100011011000;
    assign parity_check_matrix[1809] = 12'b011100100111;
    assign parity_check_matrix[1810] = 12'b001101011000;
    assign parity_check_matrix[1811] = 12'b110010100111;
    assign parity_check_matrix[1812] = 12'b010101011000;
    assign parity_check_matrix[1813] = 12'b101010100111;
    assign parity_check_matrix[1814] = 12'b100101011000;
    assign parity_check_matrix[1815] = 12'b011010100111;
    assign parity_check_matrix[1816] = 12'b011001011000;
    assign parity_check_matrix[1817] = 12'b100110100111;
    assign parity_check_matrix[1818] = 12'b101001011000;
    assign parity_check_matrix[1819] = 12'b010110100111;
    assign parity_check_matrix[1820] = 12'b110001011000;
    assign parity_check_matrix[1821] = 12'b001110100111;
    assign parity_check_matrix[1822] = 12'b001110011000;
    assign parity_check_matrix[1823] = 12'b110001100111;
    assign parity_check_matrix[1824] = 12'b010110011000;
    assign parity_check_matrix[1825] = 12'b101001100111;
    assign parity_check_matrix[1826] = 12'b100110011000;
    assign parity_check_matrix[1827] = 12'b011001100111;
    assign parity_check_matrix[1828] = 12'b011010011000;
    assign parity_check_matrix[1829] = 12'b100101100111;
    assign parity_check_matrix[1830] = 12'b101010011000;
    assign parity_check_matrix[1831] = 12'b010101100111;
    assign parity_check_matrix[1832] = 12'b110010011000;
    assign parity_check_matrix[1833] = 12'b001101100111;
    assign parity_check_matrix[1834] = 12'b011100011000;
    assign parity_check_matrix[1835] = 12'b100011100111;
    assign parity_check_matrix[1836] = 12'b101100011000;
    assign parity_check_matrix[1837] = 12'b010011100111;
    assign parity_check_matrix[1838] = 12'b110100011000;
    assign parity_check_matrix[1839] = 12'b001011100111;
    assign parity_check_matrix[1840] = 12'b111000011000;
    assign parity_check_matrix[1841] = 12'b000111100111;
    assign parity_check_matrix[1842] = 12'b000111101000;
    assign parity_check_matrix[1843] = 12'b111000010111;
    assign parity_check_matrix[1844] = 12'b001011101000;
    assign parity_check_matrix[1845] = 12'b110100010111;
    assign parity_check_matrix[1846] = 12'b010011101000;
    assign parity_check_matrix[1847] = 12'b101100010111;
    assign parity_check_matrix[1848] = 12'b100011101000;
    assign parity_check_matrix[1849] = 12'b011100010111;
    assign parity_check_matrix[1850] = 12'b001101101000;
    assign parity_check_matrix[1851] = 12'b110010010111;
    assign parity_check_matrix[1852] = 12'b010101101000;
    assign parity_check_matrix[1853] = 12'b101010010111;
    assign parity_check_matrix[1854] = 12'b100101101000;
    assign parity_check_matrix[1855] = 12'b011010010111;
    assign parity_check_matrix[1856] = 12'b011001101000;
    assign parity_check_matrix[1857] = 12'b100110010111;
    assign parity_check_matrix[1858] = 12'b101001101000;
    assign parity_check_matrix[1859] = 12'b010110010111;
    assign parity_check_matrix[1860] = 12'b110001101000;
    assign parity_check_matrix[1861] = 12'b001110010111;
    assign parity_check_matrix[1862] = 12'b001110101000;
    assign parity_check_matrix[1863] = 12'b110001010111;
    assign parity_check_matrix[1864] = 12'b010110101000;
    assign parity_check_matrix[1865] = 12'b101001010111;
    assign parity_check_matrix[1866] = 12'b100110101000;
    assign parity_check_matrix[1867] = 12'b011001010111;
    assign parity_check_matrix[1868] = 12'b011010101000;
    assign parity_check_matrix[1869] = 12'b100101010111;
    assign parity_check_matrix[1870] = 12'b101010101000;
    assign parity_check_matrix[1871] = 12'b010101010111;
    assign parity_check_matrix[1872] = 12'b110010101000;
    assign parity_check_matrix[1873] = 12'b001101010111;
    assign parity_check_matrix[1874] = 12'b011100101000;
    assign parity_check_matrix[1875] = 12'b100011010111;
    assign parity_check_matrix[1876] = 12'b101100101000;
    assign parity_check_matrix[1877] = 12'b010011010111;
    assign parity_check_matrix[1878] = 12'b110100101000;
    assign parity_check_matrix[1879] = 12'b001011010111;
    assign parity_check_matrix[1880] = 12'b111000101000;
    assign parity_check_matrix[1881] = 12'b000111010111;
    assign parity_check_matrix[1882] = 12'b001111001000;
    assign parity_check_matrix[1883] = 12'b110000110111;
    assign parity_check_matrix[1884] = 12'b010111001000;
    assign parity_check_matrix[1885] = 12'b101000110111;
    assign parity_check_matrix[1886] = 12'b100111001000;
    assign parity_check_matrix[1887] = 12'b011000110111;
    assign parity_check_matrix[1888] = 12'b011011001000;
    assign parity_check_matrix[1889] = 12'b100100110111;
    assign parity_check_matrix[1890] = 12'b101011001000;
    assign parity_check_matrix[1891] = 12'b010100110111;
    assign parity_check_matrix[1892] = 12'b110011001000;
    assign parity_check_matrix[1893] = 12'b001100110111;
    assign parity_check_matrix[1894] = 12'b011101001000;
    assign parity_check_matrix[1895] = 12'b100010110111;
    assign parity_check_matrix[1896] = 12'b101101001000;
    assign parity_check_matrix[1897] = 12'b010010110111;
    assign parity_check_matrix[1898] = 12'b110101001000;
    assign parity_check_matrix[1899] = 12'b001010110111;
    assign parity_check_matrix[1900] = 12'b111001001000;
    assign parity_check_matrix[1901] = 12'b000110110111;
    assign parity_check_matrix[1902] = 12'b011110001000;
    assign parity_check_matrix[1903] = 12'b100001110111;
    assign parity_check_matrix[1904] = 12'b101110001000;
    assign parity_check_matrix[1905] = 12'b010001110111;
    assign parity_check_matrix[1906] = 12'b110110001000;
    assign parity_check_matrix[1907] = 12'b001001110111;
    assign parity_check_matrix[1908] = 12'b111010001000;
    assign parity_check_matrix[1909] = 12'b000101110111;
    assign parity_check_matrix[1910] = 12'b111100001000;
    assign parity_check_matrix[1911] = 12'b000011110111;
    assign parity_check_matrix[1912] = 12'b000111110000;
    assign parity_check_matrix[1913] = 12'b111000001111;
    assign parity_check_matrix[1914] = 12'b001011110000;
    assign parity_check_matrix[1915] = 12'b110100001111;
    assign parity_check_matrix[1916] = 12'b010011110000;
    assign parity_check_matrix[1917] = 12'b101100001111;
    assign parity_check_matrix[1918] = 12'b100011110000;
    assign parity_check_matrix[1919] = 12'b011100001111;
    assign parity_check_matrix[1920] = 12'b001101110000;
    assign parity_check_matrix[1921] = 12'b110010001111;
    assign parity_check_matrix[1922] = 12'b010101110000;
    assign parity_check_matrix[1923] = 12'b101010001111;
    assign parity_check_matrix[1924] = 12'b100101110000;
    assign parity_check_matrix[1925] = 12'b011010001111;
    assign parity_check_matrix[1926] = 12'b011001110000;
    assign parity_check_matrix[1927] = 12'b100110001111;
    assign parity_check_matrix[1928] = 12'b101001110000;
    assign parity_check_matrix[1929] = 12'b010110001111;
    assign parity_check_matrix[1930] = 12'b110001110000;
    assign parity_check_matrix[1931] = 12'b001110001111;
    assign parity_check_matrix[1932] = 12'b001110110000;
    assign parity_check_matrix[1933] = 12'b110001001111;
    assign parity_check_matrix[1934] = 12'b010110110000;
    assign parity_check_matrix[1935] = 12'b101001001111;
    assign parity_check_matrix[1936] = 12'b100110110000;
    assign parity_check_matrix[1937] = 12'b011001001111;
    assign parity_check_matrix[1938] = 12'b011010110000;
    assign parity_check_matrix[1939] = 12'b100101001111;
    assign parity_check_matrix[1940] = 12'b101010110000;
    assign parity_check_matrix[1941] = 12'b010101001111;
    assign parity_check_matrix[1942] = 12'b110010110000;
    assign parity_check_matrix[1943] = 12'b001101001111;
    assign parity_check_matrix[1944] = 12'b011100110000;
    assign parity_check_matrix[1945] = 12'b100011001111;
    assign parity_check_matrix[1946] = 12'b101100110000;
    assign parity_check_matrix[1947] = 12'b010011001111;
    assign parity_check_matrix[1948] = 12'b110100110000;
    assign parity_check_matrix[1949] = 12'b001011001111;
    assign parity_check_matrix[1950] = 12'b111000110000;
    assign parity_check_matrix[1951] = 12'b000111001111;
    assign parity_check_matrix[1952] = 12'b001111010000;
    assign parity_check_matrix[1953] = 12'b110000101111;
    assign parity_check_matrix[1954] = 12'b010111010000;
    assign parity_check_matrix[1955] = 12'b101000101111;
    assign parity_check_matrix[1956] = 12'b100111010000;
    assign parity_check_matrix[1957] = 12'b011000101111;
    assign parity_check_matrix[1958] = 12'b011011010000;
    assign parity_check_matrix[1959] = 12'b100100101111;
    assign parity_check_matrix[1960] = 12'b101011010000;
    assign parity_check_matrix[1961] = 12'b010100101111;
    assign parity_check_matrix[1962] = 12'b110011010000;
    assign parity_check_matrix[1963] = 12'b001100101111;
    assign parity_check_matrix[1964] = 12'b011101010000;
    assign parity_check_matrix[1965] = 12'b100010101111;
    assign parity_check_matrix[1966] = 12'b101101010000;
    assign parity_check_matrix[1967] = 12'b010010101111;
    assign parity_check_matrix[1968] = 12'b110101010000;
    assign parity_check_matrix[1969] = 12'b001010101111;
    assign parity_check_matrix[1970] = 12'b111001010000;
    assign parity_check_matrix[1971] = 12'b000110101111;
    assign parity_check_matrix[1972] = 12'b011110010000;
    assign parity_check_matrix[1973] = 12'b100001101111;
    assign parity_check_matrix[1974] = 12'b101110010000;
    assign parity_check_matrix[1975] = 12'b010001101111;
    assign parity_check_matrix[1976] = 12'b110110010000;
    assign parity_check_matrix[1977] = 12'b001001101111;
    assign parity_check_matrix[1978] = 12'b111010010000;
    assign parity_check_matrix[1979] = 12'b000101101111;
    assign parity_check_matrix[1980] = 12'b111100010000;
    assign parity_check_matrix[1981] = 12'b000011101111;
    assign parity_check_matrix[1982] = 12'b001111100000;
    assign parity_check_matrix[1983] = 12'b110000011111;
    assign parity_check_matrix[1984] = 12'b010111100000;
    assign parity_check_matrix[1985] = 12'b101000011111;
    assign parity_check_matrix[1986] = 12'b100111100000;
    assign parity_check_matrix[1987] = 12'b011000011111;
    assign parity_check_matrix[1988] = 12'b011011100000;
    assign parity_check_matrix[1989] = 12'b100100011111;
    assign parity_check_matrix[1990] = 12'b101011100000;
    assign parity_check_matrix[1991] = 12'b010100011111;
    assign parity_check_matrix[1992] = 12'b110011100000;
    assign parity_check_matrix[1993] = 12'b001100011111;
    assign parity_check_matrix[1994] = 12'b011101100000;
    assign parity_check_matrix[1995] = 12'b100010011111;
    assign parity_check_matrix[1996] = 12'b101101100000;
    assign parity_check_matrix[1997] = 12'b010010011111;
    assign parity_check_matrix[1998] = 12'b110101100000;
    assign parity_check_matrix[1999] = 12'b001010011111;
    assign parity_check_matrix[2000] = 12'b111001100000;
    assign parity_check_matrix[2001] = 12'b000110011111;
    assign parity_check_matrix[2002] = 12'b011110100000;
    assign parity_check_matrix[2003] = 12'b100001011111;
    assign parity_check_matrix[2004] = 12'b101110100000;
    assign parity_check_matrix[2005] = 12'b010001011111;
    assign parity_check_matrix[2006] = 12'b110110100000;
    assign parity_check_matrix[2007] = 12'b001001011111;
    assign parity_check_matrix[2008] = 12'b111010100000;
    assign parity_check_matrix[2009] = 12'b000101011111;
    assign parity_check_matrix[2010] = 12'b111100100000;
    assign parity_check_matrix[2011] = 12'b000011011111;
    assign parity_check_matrix[2012] = 12'b011111000000;
    assign parity_check_matrix[2013] = 12'b100000111111;
    assign parity_check_matrix[2014] = 12'b101111000000;
    assign parity_check_matrix[2015] = 12'b010000111111;
    assign parity_check_matrix[2016] = 12'b110111000000;
    assign parity_check_matrix[2017] = 12'b001000111111;
    assign parity_check_matrix[2018] = 12'b111011000000;
    assign parity_check_matrix[2019] = 12'b000100111111;
    assign parity_check_matrix[2020] = 12'b111101000000;
    assign parity_check_matrix[2021] = 12'b000010111111;
    assign parity_check_matrix[2022] = 12'b111110000000;
    assign parity_check_matrix[2023] = 12'b000001111111;
    assign parity_check_matrix[2024] = 12'b011111111111;
    assign parity_check_matrix[2025] = 12'b101111111111;
    assign parity_check_matrix[2026] = 12'b110111111111;
    assign parity_check_matrix[2027] = 12'b111011111111;
    assign parity_check_matrix[2028] = 12'b111101111111;
    assign parity_check_matrix[2029] = 12'b111110111111;
    assign parity_check_matrix[2030] = 12'b111111011111;
    assign parity_check_matrix[2031] = 12'b111111101111;
    assign parity_check_matrix[2032] = 12'b111111110111;
    assign parity_check_matrix[2033] = 12'b111111111011;
    assign parity_check_matrix[2034] = 12'b111111111101;
    assign parity_check_matrix[2035] = 12'b111111111110;
    assign parity_check_matrix[2036] = 12'b100000000000;
    assign parity_check_matrix[2037] = 12'b010000000000;
    assign parity_check_matrix[2038] = 12'b001000000000;
    assign parity_check_matrix[2039] = 12'b000100000000;
    assign parity_check_matrix[2040] = 12'b000010000000;
    assign parity_check_matrix[2041] = 12'b000001000000;
    assign parity_check_matrix[2042] = 12'b000000100000;
    assign parity_check_matrix[2043] = 12'b000000010000;
    assign parity_check_matrix[2044] = 12'b000000001000;
    assign parity_check_matrix[2045] = 12'b000000000100;
    assign parity_check_matrix[2046] = 12'b000000000010;
    assign parity_check_matrix[2047] = 12'b000000000001;
  end else begin : gen_default_parity
    `BR_ASSERT_STATIC(invalid_parity_width_a, 1'b0)
  end

  // ri lint_check_on EXPR_ID_LIMIT

  //------
  // Optionally register the syndrome before decoding.
  //------
  logic internal_valid;
  logic [CodewordWidth-1:0] internal_codeword;
  logic [ParityWidth-1:0] internal_error_syndrome;

  br_delay_valid #(
      .Width(CodewordWidth + ParityWidth),
      .NumStages(RegisterSyndrome),
      .EnableAssertFinalNotValid(EnableAssertFinalNotValid)
  ) br_delay_valid_syndrome (
      .clk,
      .rst,
      .in_valid(rcv_valid_d),
      .in({cw, syndrome}),
      .out_valid(internal_valid),
      .out({internal_codeword, internal_error_syndrome}),
      .out_valid_stages(),  // unused
      .out_stages()  // unused
  );

  //------
  // Decode syndrome.
  //------
  // * Case 0: Syndrome is zero, no errors detected.
  // * Case 1: Syndrome is for a nonzero even number of bits in error, which happens when
  //   the syndrome is nonzero and even in a Hsiao SECDED code.
  //   Maximum likelihood decoding produces multiple equiprobable candidate codewords, so
  //   treat as detected-but-uncorrectable.
  //   NOTE: We are returning *some* message but it is likely to have been corrupted!
  // * Case 2: Syndrome is for an odd number of bits in error, which happens when the syndrome
  //   is odd in a Hsiao SECDED code.
  //   * Case 2a: Rarely this can be a three-bit error that is actually detected-but-uncorrectable.
  //   * Case 2b: Usually this is a single-bit error, which is always closest to exactly one codeword.
  //     So with maximum likelihood decoding we can correct it.
  logic internal_error_syndrome_parity;
  logic internal_error_syndrome_is_zero;
  logic internal_error_syndrome_is_even;
  logic internal_error_syndrome_is_odd;

  assign internal_error_syndrome_parity  = ^internal_error_syndrome;
  assign internal_error_syndrome_is_zero = internal_error_syndrome == '0;
  assign internal_error_syndrome_is_even = !internal_error_syndrome_parity;
  assign internal_error_syndrome_is_odd  = internal_error_syndrome_parity;

  // Case 0 (no errors detected) -- implicitly true if case 1, 2a, and 2b are all false.

  // Case 1 (detected-but-uncorrectable with nonzero and even syndrome)
  logic internal_due_even;
  assign internal_due_even = !internal_error_syndrome_is_zero && internal_error_syndrome_is_even;

  // Case 2 - need more information to decide if it's case 2a or 2b.
  logic [CodewordWidth-1:0] internal_h_column_match;
  for (genvar i = 0; i < CodewordWidth; i++) begin : gen_col_match
    assign internal_h_column_match[i] = (internal_error_syndrome == parity_check_matrix[i]);
  end

  // Case 2a (detected-but-uncorrectable with odd syndrome)
  // This happens when the syndrome is odd but it doesn't match any of the columns in H.
  // Since the code is guaranteed to correct any single-bit error, this means it must be
  // an odd number (at least 3) of bits in error.
  logic internal_due_odd;
  assign internal_due_odd = internal_error_syndrome_is_odd && (internal_h_column_match == '0);

  // Merge case 1 and 2a (detected-but-uncorrectable)
  logic internal_error_due;
  assign internal_error_due = (internal_due_even || internal_due_odd);

  // Case 2b (correctable with single-bit error)
  logic internal_error_ce;
  assign internal_error_ce =
    internal_error_syndrome_is_odd && (internal_h_column_match != '0);

  //------
  // Correct the codeword (if necessary and possible), then extract the message and data.
  //------
  // If there was a DUE, then the corr codeword is still corrupted and
  // the message and data are likely to also be corrupted.

  logic [CodewordWidth-1:0] internal_corrected_codeword;

  assign internal_corrected_codeword = internal_codeword ^ internal_h_column_match;

  `BR_ASSERT_IMPL(internal_h_column_match_onehot0_a,
                  internal_valid |-> $onehot0(internal_h_column_match))
  `BR_ASSERT_IMPL(due_no_h_column_match_a,
                  internal_valid && internal_error_due |->
                  (internal_h_column_match == '0))
  `BR_ASSERT_IMPL(no_error_correction_a,
                  internal_valid && !internal_error_ce |->
                  (internal_corrected_codeword == internal_codeword))
  `BR_ASSERT_IMPL(error_correction_a,
                  internal_valid && internal_error_ce |->
                  (internal_corrected_codeword != internal_codeword))

  //------
  // Optionally register the output signals.
  //------
  logic [InputWidth-1:0] internal_corrected_codeword_compressed;
  assign `BR_INSERT_TO_MSB(internal_corrected_codeword_compressed, internal_corrected_codeword[CodewordWidth-1 -: ParityWidth])
  assign `BR_INSERT_TO_LSB(internal_corrected_codeword_compressed, internal_corrected_codeword[DataWidth-1:0])
  if (CodewordWidth > InputWidth) begin : gen_internal_corrected_codeword_unused
    `BR_UNUSED_NAMED(unused_internal_corrected_codeword, internal_corrected_codeword[MessageWidth-1 : DataWidth])
  end
  br_delay_valid #(
      .Width(InputWidth + 2 + ParityWidth),
      .NumStages(RegisterOutputs == 1 ? 1 : 0),
      .EnableAssertFinalNotValid(EnableAssertFinalNotValid)
  ) br_delay_valid_outputs (
      .clk,
      .rst,
      .in_valid(internal_valid),
      .in({internal_corrected_codeword_compressed,
          internal_error_ce,
          internal_error_due,
          internal_error_syndrome}),
      .out_valid(dec_valid),
      .out({dec_codeword,
            dec_error_ce,
            dec_error_due,
            dec_error_syndrome}),
      .out_valid_stages(),  // unused
      .out_stages()  // unused
  );

  // ri lint_check_waive FULL_RANGE
  assign dec_data = dec_codeword[DataWidth-1:0];

  //------------------------------------------
  // Implementation checks
  //------------------------------------------
  `BR_ASSERT_IMPL(latency_a, rcv_valid |-> ##Latency dec_valid)
  `BR_ASSERT_IMPL(ce_due_mutually_exclusive_a,
                  dec_valid |-> $onehot0({dec_error_ce, dec_error_due}))
  `BR_COVER_IMPL(ce_c, dec_valid && dec_error_ce)
  `BR_COVER_IMPL(due_c, dec_valid && dec_error_due)

  // verilog_format: on
  // verilog_lint: waive-stop line-length

endmodule : br_ecc_secded_decoder
