// SPDX-License-Identifier: Apache-2.0

`include "br_asserts_internal.svh"

module br_fifo_shared_pstatic_ctrl #(
    // Number of logical FIFOs. Must be >=2.
    parameter int NumFifos = 2,
    // Total depth of the FIFO.
    // Must be greater than or equal to the number of logical FIFOs.
    parameter int Depth = 2,
    // Width of the data. Must be >=1.
    parameter int Width = 1,
    // The depth of the pop-side staging buffer.
    // This affects the pop bandwidth of each logical FIFO.
    // The bandwidth will be `StagingBufferDepth / (PointerRamReadLatency + 1)`.
    parameter int StagingBufferDepth = 1,
    // If 1, make sure pop_valid/pop_data are registered at the output
    // of the staging buffer. This adds a cycle of cut-through latency.
    parameter bit RegisterPopOutputs = 0,
    // The number of cycles between ram read address and read data. Must be >=0.
    parameter int RamReadLatency = 0,
    // If 1, cover that the push side experiences backpressure.
    // If 0, assert that there is never backpressure.
    parameter bit EnableCoverPushBackpressure = 1,
    // If 1, assert that push_valid is stable when backpressured.
    // If 0, cover that push_valid can be unstable.
    parameter bit EnableAssertPushValidStability = EnableCoverPushBackpressure,
    // If 1, assert that push_data is stable when backpressured.
    // If 0, cover that push_data can be unstable.
    // ri lint_check_waive PARAM_NOT_USED
    parameter bit EnableAssertPushDataStability = EnableAssertPushValidStability,
    // If 1, assert that push_data is always known (not X) when push_valid is asserted.
    parameter bit EnableAssertPushDataKnown = 1,
    // If 1, then assert there are no valid bits asserted and that the FIFO is
    // empty at the end of the test.
    // ri lint_check_waive PARAM_NOT_USED
    parameter bit EnableAssertFinalNotValid = 1,

    localparam int FifoIdWidth = br_math::clamped_clog2(NumFifos),
    localparam int AddrWidth   = br_math::clamped_clog2(Depth),
    localparam int CountWidth  = $clog2(Depth + 1)
) (
    input logic clk,
    input logic rst,

    // Fifo configuration
    // These can come from straps or CSRs, but they must be set before reset is
    // deasserted and then held stable until reset is asserted.
    // The base and bound addresses determine the range of RAM addresses given
    // to each logical FIFO. They are both inclusive, so logical FIFO i will
    // increment from config_base[i] up to config_bound[i] before wrapping back
    // around to config_base[i] again.
    // The minimum size for a given logical FIFO is 1, meaning that
    // config_bound[i] must be >= config_base[i] for all i.
    // The address ranges must be in ascending order.
    input logic [NumFifos-1:0][AddrWidth-1:0] config_base,
    input logic [NumFifos-1:0][AddrWidth-1:0] config_bound,
    // Error is asserted if the base and bound addresses are misconfigured.
    // For instance, if any address is >= Depth, config_base[i] > config_bound[i],
    // or config_base[i] <= config_bound[i-1] for i > 0.
    output logic config_error,

    // Push-side interface
    output logic                   push_ready,
    input  logic                   push_valid,
    input  logic [      Width-1:0] push_data,
    input  logic [FifoIdWidth-1:0] push_fifo_id,
    output logic [   NumFifos-1:0] push_full,

    // Pop-side interface
    input  logic [NumFifos-1:0]            pop_ready,
    output logic [NumFifos-1:0]            pop_valid,
    output logic [NumFifos-1:0][Width-1:0] pop_data,
    output logic [NumFifos-1:0]            pop_empty,

    // RAM read/write ports
    output logic                 ram_wr_valid,
    output logic [AddrWidth-1:0] ram_wr_addr,
    output logic [    Width-1:0] ram_wr_data,
    output logic                 ram_rd_addr_valid,
    output logic [AddrWidth-1:0] ram_rd_addr,
    input  logic                 ram_rd_data_valid,
    input  logic [    Width-1:0] ram_rd_data
);

  // Integration assertions
  `BR_ASSERT_STATIC(num_fifos_gte_2_a, NumFifos >= 2)
  `BR_ASSERT_STATIC(depth_gte_num_fifos_a, Depth >= NumFifos)
  `BR_ASSERT_STATIC(width_gte_1_a, Width >= 1)

  // Other integration checks in submodules

  // Implementation
  logic [NumFifos-1:0][CountWidth-1:0] config_size;

  br_fifo_shared_pstatic_size_calc #(
      .NumFifos(NumFifos),
      .Depth(Depth)
  ) br_fifo_shared_pstatic_size_calc (
      .clk,
      .rst,
      .config_base,
      .config_bound,
      .config_size,
      .config_error
  );

  logic [NumFifos-1:0] advance_tail;
  logic [NumFifos-1:0][AddrWidth-1:0] tail_next;
  logic [NumFifos-1:0][AddrWidth-1:0] tail;

  br_fifo_shared_pstatic_push_ctrl #(
      .NumFifos(NumFifos),
      .Depth(Depth),
      .Width(Width),
      .EnableCoverPushBackpressure(EnableCoverPushBackpressure),
      .EnableAssertPushValidStability(EnableAssertPushValidStability),
      .EnableAssertPushDataStability(EnableAssertPushDataStability),
      .EnableAssertPushDataKnown(EnableAssertPushDataKnown),
      .EnableAssertFinalNotValid(EnableAssertFinalNotValid)
  ) br_fifo_shared_pstatic_push_ctrl (
      .clk,
      .rst,
      .config_base,
      .config_bound,
      .push_ready,
      .push_valid,
      .push_data,
      .push_fifo_id,
      .push_full,
      .ram_wr_valid,
      .ram_wr_addr,
      .ram_wr_data,
      .advance_tail,
      .tail_next,
      .tail
  );

  logic [NumFifos-1:0] head_ready;
  logic [NumFifos-1:0] head_valid;
  logic [NumFifos-1:0][AddrWidth-1:0] head;
  logic [NumFifos-1:0] ram_empty;
  logic [NumFifos-1:0][CountWidth-1:0] ram_items;

  br_fifo_shared_pstatic_ptr_mgr #(
      .NumFifos(NumFifos),
      .Depth(Depth),
      // Keep this at 0 for now to avoid introducing extra registers.
      // May expose this as a top-level parameter if there is a timing issue.
      .RegisterRamItems(0),
      .EnableAssertFinalNotValid(EnableAssertFinalNotValid)
  ) br_fifo_shared_pstatic_ptr_mgr (
      .clk,
      .rst,
      .config_base,
      .config_bound,
      .config_size,
      .advance_tail,
      .tail_next,
      .tail,
      .push_full,
      .head_ready,
      .head_valid,
      .head,
      .ram_empty,
      .ram_items
  );

  br_fifo_shared_pop_ctrl #(
      .NumReadPorts(1),
      .NumFifos(NumFifos),
      .Depth(Depth),
      .Width(Width),
      .StagingBufferDepth(StagingBufferDepth),
      .RegisterPopOutputs(RegisterPopOutputs),
      .RamReadLatency(RamReadLatency)
  ) br_fifo_shared_pop_ctrl (
      .clk,
      .rst,
      .head_valid,
      .head_ready,
      .head,
      .ram_empty,
      .ram_items,
      .pop_valid,
      .pop_ready,
      .pop_data,
      .pop_empty,
      .dealloc_valid(),  // Not used
      .dealloc_entry_id(),  // Not used
      .data_ram_rd_addr_valid(ram_rd_addr_valid),
      .data_ram_rd_addr(ram_rd_addr),
      .data_ram_rd_data_valid(ram_rd_data_valid),
      .data_ram_rd_data(ram_rd_data)
  );
endmodule
