// Copyright 2024 The Bedrock-RTL Authors
//
// Licensed under the Apache License, Version 2.0 (the "License");
// Copyright 2024 The Bedrock-RTL Authors
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//     http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.

// Bedrock-RTL Single-Error-Correcting, Double-Error-Detecting (SECDED - Hsiao) Decoder
//
// Decodes a codeword using a single-error-correcting, double-error-detecting
// linear block code in systematic form (in layperson's terms: a Hsiao SECDED [1] decoder,
// closely related to Hamming codes).
//
// Systematic form means that the codeword is formed by appending the
// calculated parity bits to the message, i.e., the code has the property
// that the message bits are 1:1 with a slice of bits in the codeword (if they
// have not been corrupted).
//
// In Bedrock ECC libs, our convention is to always append the parity bits on
// the MSbs:
//     codeword == {parity, message}
//
// This is a purely combinational module. Valid bits are provided for
// convenience of user integration and port compatibility with the
// corresponding encoder module (br_ecc_secded_encoder).
//
// The data is still marked valid even if an error is detected.
//
// Any data width >= 1 is supported. It is considered internally zero-padded up to
// the nearest power-of-2 message width as part of decoding. The following
// table outlines the number of parity bits required for different message widths.
//
// | Message Width (k) | Parity Width (r) | Codeword Width (n)|
// |-------------------|------------------|-------------------|
// | 4                 | 4                | 8                 |
// | 8                 | 5                | 13                |
// | 16                | 6                | 22                |
// | 32                | 7                | 39                |
// | 64                | 8                | 72                |
// | 128               | 9                | 137               |
// | 256               | 10               | 266               |
// | 512               | 11               | 523               |
// | 1024              | 12               | 1036              |
//
// The number of parity bits must be one of the values in the table above
// or the module will not elaborate.
//
// References:
// [1] https://ieeexplore.ieee.org/abstract/document/5391627

`include "br_asserts_internal.svh"

// TODO(mgottscho): Pipeline the syndrome decoding and then correction with a parameter.
module br_ecc_secded_decoder #(
    parameter int DataWidth = 1,  // Must be at least 1
    parameter int ParityWidth = 4,  // Must be at least 4 and at most 12
    localparam int MessageWidth = 2 ** $clog2(DataWidth),
    localparam int CodewordWidth = MessageWidth + ParityWidth
) (
    input  logic                     codeword_valid,
    input  logic [CodewordWidth-1:0] codeword,
    output logic                     data_valid,
    output logic [    DataWidth-1:0] data,
    output logic                     error_valid,
    output logic                     error_corrected,
    output logic                     error_detected_but_uncorrectable,
    output logic [  ParityWidth-1:0] error_syndrome
);

  //------------------------------------------
  // Integration checks
  //------------------------------------------
  `BR_ASSERT_STATIC(message_width_gte_1_a, DataWidth >= 1)
  `BR_ASSERT_STATIC(parity_width_gte_4_a, ParityWidth >= 4)
  `BR_ASSERT_STATIC(parity_width_lte_12_a, ParityWidth <= 12)
  `BR_ASSERT_STATIC(message_width_is_power_of_2_a, br_math::is_power_of_2(MessageWidth))

  //------------------------------------------
  // Implementation
  //------------------------------------------

  // verilog_format: off
  // verilog_lint: waive-start line-length
  if (CodewordWidth == 4 && MessageWidth == 4) begin : gen_8_4
    `BR_ASSERT_STATIC(parity_width_matches_a, ParityWidth == 4)
    assign syndrome[0] = codeword[1] ^ codeword[2] ^ codeword[3] ^ codeword[4];
    assign syndrome[1] = codeword[0] ^ codeword[2] ^ codeword[3] ^ codeword[5];
    assign syndrome[2] = codeword[0] ^ codeword[1] ^ codeword[3] ^ codeword[6];
    assign syndrome[3] = codeword[0] ^ codeword[1] ^ codeword[2] ^ codeword[7];
  end else if (CodewordWidth == 13 && MessageWidth == 8) begin : gen_13_8
    `BR_ASSERT_STATIC(parity_width_matches_a, ParityWidth == 5)
    assign syndrome[0] = codeword[4] ^ codeword[5] ^ codeword[6] ^ codeword[7] ^ codeword[8];
    assign syndrome[1] = codeword[1] ^ codeword[2] ^ codeword[3] ^ codeword[7] ^ codeword[9];
    assign syndrome[2] = codeword[0] ^ codeword[2] ^ codeword[3] ^ codeword[5] ^ codeword[6] ^ codeword[10];
    assign syndrome[3] = codeword[0] ^ codeword[1] ^ codeword[3] ^ codeword[4] ^ codeword[6] ^ codeword[11];
    assign syndrome[4] = codeword[0] ^ codeword[1] ^ codeword[2] ^ codeword[4] ^ codeword[5] ^ codeword[7] ^ codeword[12];
  end else if (CodewordWidth == 22 && MessageWidth == 16) begin : gen_22_16
    `BR_ASSERT_STATIC(parity_width_matches_a, ParityWidth == 6)
    assign syndrome[0] = codeword[10] ^ codeword[11] ^ codeword[12] ^ codeword[13] ^ codeword[14] ^ codeword[15] ^ codeword[16];
    assign syndrome[1] = codeword[4] ^ codeword[5] ^ codeword[6] ^ codeword[7] ^ codeword[8] ^ codeword[9] ^ codeword[17];
    assign syndrome[2] = codeword[1] ^ codeword[2] ^ codeword[3] ^ codeword[7] ^ codeword[8] ^ codeword[9] ^ codeword[13] ^ codeword[14] ^ codeword[15] ^ codeword[18];
    assign syndrome[3] = codeword[0] ^ codeword[2] ^ codeword[3] ^ codeword[5] ^ codeword[6] ^ codeword[9] ^ codeword[11] ^ codeword[12] ^ codeword[15] ^ codeword[19];
    assign syndrome[4] = codeword[0] ^ codeword[1] ^ codeword[3] ^ codeword[4] ^ codeword[6] ^ codeword[8] ^ codeword[10] ^ codeword[12] ^ codeword[14] ^ codeword[20];
    assign syndrome[5] = codeword[0] ^ codeword[1] ^ codeword[2] ^ codeword[4] ^ codeword[5] ^ codeword[7] ^ codeword[10] ^ codeword[11] ^ codeword[13] ^ codeword[21];
  end else if (CodewordWidth == 39 && MessageWidth == 32) begin : gen_39_32
    `BR_ASSERT_STATIC(parity_width_matches_a, ParityWidth == 7)
    assign syndrome[0] = codeword[20] ^ codeword[21] ^ codeword[22] ^ codeword[23] ^ codeword[24] ^ codeword[25] ^ codeword[26] ^ codeword[27] ^ codeword[28] ^ codeword[29] ^ codeword[30] ^ codeword[31] ^ codeword[32];
    assign syndrome[1] = codeword[10] ^ codeword[11] ^ codeword[12] ^ codeword[13] ^ codeword[14] ^ codeword[15] ^ codeword[16] ^ codeword[17] ^ codeword[18] ^ codeword[19] ^ codeword[30] ^ codeword[31] ^ codeword[33];
    assign syndrome[2] = codeword[4] ^ codeword[5] ^ codeword[6] ^ codeword[7] ^ codeword[8] ^ codeword[9] ^ codeword[16] ^ codeword[17] ^ codeword[18] ^ codeword[19] ^ codeword[26] ^ codeword[27] ^ codeword[28] ^ codeword[29] ^ codeword[34];
    assign syndrome[3] = codeword[1] ^ codeword[2] ^ codeword[3] ^ codeword[7] ^ codeword[8] ^ codeword[9] ^ codeword[13] ^ codeword[14] ^ codeword[15] ^ codeword[19] ^ codeword[23] ^ codeword[24] ^ codeword[25] ^ codeword[29] ^ codeword[35];
    assign syndrome[4] = codeword[0] ^ codeword[2] ^ codeword[3] ^ codeword[5] ^ codeword[6] ^ codeword[9] ^ codeword[11] ^ codeword[12] ^ codeword[15] ^ codeword[18] ^ codeword[21] ^ codeword[22] ^ codeword[25] ^ codeword[28] ^ codeword[36];
    assign syndrome[5] = codeword[0] ^ codeword[1] ^ codeword[3] ^ codeword[4] ^ codeword[6] ^ codeword[8] ^ codeword[10] ^ codeword[12] ^ codeword[14] ^ codeword[17] ^ codeword[20] ^ codeword[22] ^ codeword[24] ^ codeword[27] ^ codeword[31] ^ codeword[37];
    assign syndrome[6] = codeword[0] ^ codeword[1] ^ codeword[2] ^ codeword[4] ^ codeword[5] ^ codeword[7] ^ codeword[10] ^ codeword[11] ^ codeword[13] ^ codeword[16] ^ codeword[20] ^ codeword[21] ^ codeword[23] ^ codeword[26] ^ codeword[30] ^ codeword[38];
  end else if (CodewordWidth == 72 && MessageWidth == 64) begin : gen_72_64
    `BR_ASSERT_STATIC(parity_width_matches_a, ParityWidth == 8)
    assign syndrome[0] = codeword[35] ^ codeword[36] ^ codeword[37] ^ codeword[38] ^ codeword[39] ^ codeword[40] ^ codeword[41] ^ codeword[42] ^ codeword[43] ^ codeword[44] ^ codeword[45] ^ codeword[46] ^ codeword[47] ^ codeword[48] ^ codeword[49] ^ codeword[50] ^ codeword[51] ^ codeword[52] ^ codeword[53] ^ codeword[54] ^ codeword[55] ^ codeword[64];
    assign syndrome[1] = codeword[20] ^ codeword[21] ^ codeword[22] ^ codeword[23] ^ codeword[24] ^ codeword[25] ^ codeword[26] ^ codeword[27] ^ codeword[28] ^ codeword[29] ^ codeword[30] ^ codeword[31] ^ codeword[32] ^ codeword[33] ^ codeword[34] ^ codeword[50] ^ codeword[51] ^ codeword[52] ^ codeword[53] ^ codeword[54] ^ codeword[55] ^ codeword[62] ^ codeword[63] ^ codeword[65];
    assign syndrome[2] = codeword[10] ^ codeword[11] ^ codeword[12] ^ codeword[13] ^ codeword[14] ^ codeword[15] ^ codeword[16] ^ codeword[17] ^ codeword[18] ^ codeword[19] ^ codeword[30] ^ codeword[31] ^ codeword[32] ^ codeword[33] ^ codeword[34] ^ codeword[45] ^ codeword[46] ^ codeword[47] ^ codeword[48] ^ codeword[49] ^ codeword[55] ^ codeword[57] ^ codeword[58] ^ codeword[59] ^ codeword[60] ^ codeword[61] ^ codeword[66];
    assign syndrome[3] = codeword[4] ^ codeword[5] ^ codeword[6] ^ codeword[7] ^ codeword[8] ^ codeword[9] ^ codeword[16] ^ codeword[17] ^ codeword[18] ^ codeword[19] ^ codeword[26] ^ codeword[27] ^ codeword[28] ^ codeword[29] ^ codeword[34] ^ codeword[41] ^ codeword[42] ^ codeword[43] ^ codeword[44] ^ codeword[49] ^ codeword[54] ^ codeword[56] ^ codeword[58] ^ codeword[59] ^ codeword[60] ^ codeword[61] ^ codeword[63] ^ codeword[67];
    assign syndrome[4] = codeword[1] ^ codeword[2] ^ codeword[3] ^ codeword[7] ^ codeword[8] ^ codeword[9] ^ codeword[13] ^ codeword[14] ^ codeword[15] ^ codeword[19] ^ codeword[23] ^ codeword[24] ^ codeword[25] ^ codeword[29] ^ codeword[33] ^ codeword[38] ^ codeword[39] ^ codeword[40] ^ codeword[44] ^ codeword[48] ^ codeword[53] ^ codeword[56] ^ codeword[57] ^ codeword[59] ^ codeword[60] ^ codeword[61] ^ codeword[62] ^ codeword[68];
    assign syndrome[5] = codeword[0] ^ codeword[2] ^ codeword[3] ^ codeword[5] ^ codeword[6] ^ codeword[9] ^ codeword[11] ^ codeword[12] ^ codeword[15] ^ codeword[18] ^ codeword[21] ^ codeword[22] ^ codeword[25] ^ codeword[28] ^ codeword[32] ^ codeword[36] ^ codeword[37] ^ codeword[40] ^ codeword[43] ^ codeword[47] ^ codeword[52] ^ codeword[56] ^ codeword[57] ^ codeword[58] ^ codeword[60] ^ codeword[61] ^ codeword[62] ^ codeword[63] ^ codeword[69];
    assign syndrome[6] = codeword[0] ^ codeword[1] ^ codeword[3] ^ codeword[4] ^ codeword[6] ^ codeword[8] ^ codeword[10] ^ codeword[12] ^ codeword[14] ^ codeword[17] ^ codeword[20] ^ codeword[22] ^ codeword[24] ^ codeword[27] ^ codeword[31] ^ codeword[35] ^ codeword[37] ^ codeword[39] ^ codeword[42] ^ codeword[46] ^ codeword[51] ^ codeword[56] ^ codeword[57] ^ codeword[58] ^ codeword[59] ^ codeword[61] ^ codeword[62] ^ codeword[63] ^ codeword[70];
    assign syndrome[7] = codeword[0] ^ codeword[1] ^ codeword[2] ^ codeword[4] ^ codeword[5] ^ codeword[7] ^ codeword[10] ^ codeword[11] ^ codeword[13] ^ codeword[16] ^ codeword[20] ^ codeword[21] ^ codeword[23] ^ codeword[26] ^ codeword[30] ^ codeword[35] ^ codeword[36] ^ codeword[38] ^ codeword[41] ^ codeword[45] ^ codeword[50] ^ codeword[56] ^ codeword[57] ^ codeword[58] ^ codeword[59] ^ codeword[60] ^ codeword[62] ^ codeword[63] ^ codeword[71];
  end else if (CodewordWidth == 137 && MessageWidth == 128) begin : gen_137_128
    `BR_ASSERT_STATIC(parity_width_matches_a, ParityWidth == 9)
    assign syndrome[0] = codeword[56] ^ codeword[57] ^ codeword[58] ^ codeword[59] ^ codeword[60] ^ codeword[61] ^ codeword[62] ^ codeword[63] ^ codeword[64] ^ codeword[65] ^ codeword[66] ^ codeword[67] ^ codeword[68] ^ codeword[69] ^ codeword[70] ^ codeword[71] ^ codeword[72] ^ codeword[73] ^ codeword[74] ^ codeword[75] ^ codeword[76] ^ codeword[77] ^ codeword[78] ^ codeword[79] ^ codeword[80] ^ codeword[81] ^ codeword[82] ^ codeword[83] ^ codeword[128];
    assign syndrome[1] = codeword[35] ^ codeword[36] ^ codeword[37] ^ codeword[38] ^ codeword[39] ^ codeword[40] ^ codeword[41] ^ codeword[42] ^ codeword[43] ^ codeword[44] ^ codeword[45] ^ codeword[46] ^ codeword[47] ^ codeword[48] ^ codeword[49] ^ codeword[50] ^ codeword[51] ^ codeword[52] ^ codeword[53] ^ codeword[54] ^ codeword[55] ^ codeword[77] ^ codeword[78] ^ codeword[79] ^ codeword[80] ^ codeword[81] ^ codeword[82] ^ codeword[83] ^ codeword[105] ^ codeword[106] ^ codeword[107] ^ codeword[108] ^ codeword[109] ^ codeword[110] ^ codeword[111] ^ codeword[112] ^ codeword[113] ^ codeword[114] ^ codeword[115] ^ codeword[116] ^ codeword[117] ^ codeword[118] ^ codeword[119] ^ codeword[120] ^ codeword[121] ^ codeword[122] ^ codeword[123] ^ codeword[124] ^ codeword[125] ^ codeword[126] ^ codeword[127] ^ codeword[129];
    assign syndrome[2] = codeword[20] ^ codeword[21] ^ codeword[22] ^ codeword[23] ^ codeword[24] ^ codeword[25] ^ codeword[26] ^ codeword[27] ^ codeword[28] ^ codeword[29] ^ codeword[30] ^ codeword[31] ^ codeword[32] ^ codeword[33] ^ codeword[34] ^ codeword[50] ^ codeword[51] ^ codeword[52] ^ codeword[53] ^ codeword[54] ^ codeword[55] ^ codeword[71] ^ codeword[72] ^ codeword[73] ^ codeword[74] ^ codeword[75] ^ codeword[76] ^ codeword[83] ^ codeword[90] ^ codeword[91] ^ codeword[92] ^ codeword[93] ^ codeword[94] ^ codeword[95] ^ codeword[96] ^ codeword[97] ^ codeword[98] ^ codeword[99] ^ codeword[100] ^ codeword[101] ^ codeword[102] ^ codeword[103] ^ codeword[104] ^ codeword[120] ^ codeword[121] ^ codeword[122] ^ codeword[123] ^ codeword[124] ^ codeword[125] ^ codeword[126] ^ codeword[127] ^ codeword[130];
    assign syndrome[3] = codeword[10] ^ codeword[11] ^ codeword[12] ^ codeword[13] ^ codeword[14] ^ codeword[15] ^ codeword[16] ^ codeword[17] ^ codeword[18] ^ codeword[19] ^ codeword[30] ^ codeword[31] ^ codeword[32] ^ codeword[33] ^ codeword[34] ^ codeword[45] ^ codeword[46] ^ codeword[47] ^ codeword[48] ^ codeword[49] ^ codeword[55] ^ codeword[66] ^ codeword[67] ^ codeword[68] ^ codeword[69] ^ codeword[70] ^ codeword[76] ^ codeword[82] ^ codeword[85] ^ codeword[86] ^ codeword[87] ^ codeword[88] ^ codeword[89] ^ codeword[95] ^ codeword[96] ^ codeword[97] ^ codeword[98] ^ codeword[99] ^ codeword[100] ^ codeword[101] ^ codeword[102] ^ codeword[103] ^ codeword[104] ^ codeword[110] ^ codeword[111] ^ codeword[112] ^ codeword[113] ^ codeword[114] ^ codeword[115] ^ codeword[116] ^ codeword[117] ^ codeword[118] ^ codeword[119] ^ codeword[131];
    assign syndrome[4] = codeword[4] ^ codeword[5] ^ codeword[6] ^ codeword[7] ^ codeword[8] ^ codeword[9] ^ codeword[16] ^ codeword[17] ^ codeword[18] ^ codeword[19] ^ codeword[26] ^ codeword[27] ^ codeword[28] ^ codeword[29] ^ codeword[34] ^ codeword[41] ^ codeword[42] ^ codeword[43] ^ codeword[44] ^ codeword[49] ^ codeword[54] ^ codeword[62] ^ codeword[63] ^ codeword[64] ^ codeword[65] ^ codeword[70] ^ codeword[75] ^ codeword[81] ^ codeword[84] ^ codeword[86] ^ codeword[87] ^ codeword[88] ^ codeword[89] ^ codeword[91] ^ codeword[92] ^ codeword[93] ^ codeword[94] ^ codeword[99] ^ codeword[100] ^ codeword[101] ^ codeword[102] ^ codeword[103] ^ codeword[104] ^ codeword[106] ^ codeword[107] ^ codeword[108] ^ codeword[109] ^ codeword[114] ^ codeword[115] ^ codeword[116] ^ codeword[117] ^ codeword[118] ^ codeword[119] ^ codeword[124] ^ codeword[125] ^ codeword[126] ^ codeword[127] ^ codeword[132];
    assign syndrome[5] = codeword[1] ^ codeword[2] ^ codeword[3] ^ codeword[7] ^ codeword[8] ^ codeword[9] ^ codeword[13] ^ codeword[14] ^ codeword[15] ^ codeword[19] ^ codeword[23] ^ codeword[24] ^ codeword[25] ^ codeword[29] ^ codeword[33] ^ codeword[38] ^ codeword[39] ^ codeword[40] ^ codeword[44] ^ codeword[48] ^ codeword[53] ^ codeword[59] ^ codeword[60] ^ codeword[61] ^ codeword[65] ^ codeword[69] ^ codeword[74] ^ codeword[80] ^ codeword[84] ^ codeword[85] ^ codeword[87] ^ codeword[88] ^ codeword[89] ^ codeword[90] ^ codeword[92] ^ codeword[93] ^ codeword[94] ^ codeword[96] ^ codeword[97] ^ codeword[98] ^ codeword[102] ^ codeword[103] ^ codeword[104] ^ codeword[105] ^ codeword[107] ^ codeword[108] ^ codeword[109] ^ codeword[111] ^ codeword[112] ^ codeword[113] ^ codeword[117] ^ codeword[118] ^ codeword[119] ^ codeword[121] ^ codeword[122] ^ codeword[123] ^ codeword[127] ^ codeword[133];
    assign syndrome[6] = codeword[0] ^ codeword[2] ^ codeword[3] ^ codeword[5] ^ codeword[6] ^ codeword[9] ^ codeword[11] ^ codeword[12] ^ codeword[15] ^ codeword[18] ^ codeword[21] ^ codeword[22] ^ codeword[25] ^ codeword[28] ^ codeword[32] ^ codeword[36] ^ codeword[37] ^ codeword[40] ^ codeword[43] ^ codeword[47] ^ codeword[52] ^ codeword[57] ^ codeword[58] ^ codeword[61] ^ codeword[64] ^ codeword[68] ^ codeword[73] ^ codeword[79] ^ codeword[84] ^ codeword[85] ^ codeword[86] ^ codeword[88] ^ codeword[89] ^ codeword[90] ^ codeword[91] ^ codeword[93] ^ codeword[94] ^ codeword[95] ^ codeword[97] ^ codeword[98] ^ codeword[100] ^ codeword[101] ^ codeword[104] ^ codeword[105] ^ codeword[106] ^ codeword[108] ^ codeword[109] ^ codeword[110] ^ codeword[112] ^ codeword[113] ^ codeword[115] ^ codeword[116] ^ codeword[119] ^ codeword[120] ^ codeword[122] ^ codeword[123] ^ codeword[125] ^ codeword[126] ^ codeword[134];
    assign syndrome[7] = codeword[0] ^ codeword[1] ^ codeword[3] ^ codeword[4] ^ codeword[6] ^ codeword[8] ^ codeword[10] ^ codeword[12] ^ codeword[14] ^ codeword[17] ^ codeword[20] ^ codeword[22] ^ codeword[24] ^ codeword[27] ^ codeword[31] ^ codeword[35] ^ codeword[37] ^ codeword[39] ^ codeword[42] ^ codeword[46] ^ codeword[51] ^ codeword[56] ^ codeword[58] ^ codeword[60] ^ codeword[63] ^ codeword[67] ^ codeword[72] ^ codeword[78] ^ codeword[84] ^ codeword[85] ^ codeword[86] ^ codeword[87] ^ codeword[89] ^ codeword[90] ^ codeword[91] ^ codeword[92] ^ codeword[94] ^ codeword[95] ^ codeword[96] ^ codeword[98] ^ codeword[99] ^ codeword[101] ^ codeword[103] ^ codeword[105] ^ codeword[106] ^ codeword[107] ^ codeword[109] ^ codeword[110] ^ codeword[111] ^ codeword[113] ^ codeword[114] ^ codeword[116] ^ codeword[118] ^ codeword[120] ^ codeword[121] ^ codeword[123] ^ codeword[124] ^ codeword[126] ^ codeword[135];
    assign syndrome[8] = codeword[0] ^ codeword[1] ^ codeword[2] ^ codeword[4] ^ codeword[5] ^ codeword[7] ^ codeword[10] ^ codeword[11] ^ codeword[13] ^ codeword[16] ^ codeword[20] ^ codeword[21] ^ codeword[23] ^ codeword[26] ^ codeword[30] ^ codeword[35] ^ codeword[36] ^ codeword[38] ^ codeword[41] ^ codeword[45] ^ codeword[50] ^ codeword[56] ^ codeword[57] ^ codeword[59] ^ codeword[62] ^ codeword[66] ^ codeword[71] ^ codeword[77] ^ codeword[84] ^ codeword[85] ^ codeword[86] ^ codeword[87] ^ codeword[88] ^ codeword[90] ^ codeword[91] ^ codeword[92] ^ codeword[93] ^ codeword[95] ^ codeword[96] ^ codeword[97] ^ codeword[99] ^ codeword[100] ^ codeword[102] ^ codeword[105] ^ codeword[106] ^ codeword[107] ^ codeword[108] ^ codeword[110] ^ codeword[111] ^ codeword[112] ^ codeword[114] ^ codeword[115] ^ codeword[117] ^ codeword[120] ^ codeword[121] ^ codeword[122] ^ codeword[124] ^ codeword[125] ^ codeword[127] ^ codeword[136];
  end else if (CodewordWidth == 266 && MessageWidth == 256) begin : gen_266_256
    `BR_ASSERT_STATIC(parity_width_matches_a, ParityWidth == 10)
    assign syndrome[0] = codeword[84] ^ codeword[85] ^ codeword[86] ^ codeword[87] ^ codeword[88] ^ codeword[89] ^ codeword[90] ^ codeword[91] ^ codeword[92] ^ codeword[93] ^ codeword[94] ^ codeword[95] ^ codeword[96] ^ codeword[97] ^ codeword[98] ^ codeword[99] ^ codeword[100] ^ codeword[101] ^ codeword[102] ^ codeword[103] ^ codeword[104] ^ codeword[105] ^ codeword[106] ^ codeword[107] ^ codeword[108] ^ codeword[109] ^ codeword[110] ^ codeword[111] ^ codeword[112] ^ codeword[113] ^ codeword[114] ^ codeword[115] ^ codeword[116] ^ codeword[117] ^ codeword[118] ^ codeword[119] ^ codeword[246] ^ codeword[247] ^ codeword[248] ^ codeword[249] ^ codeword[250] ^ codeword[251] ^ codeword[252] ^ codeword[253] ^ codeword[254] ^ codeword[255] ^ codeword[256];
    assign syndrome[1] = codeword[56] ^ codeword[57] ^ codeword[58] ^ codeword[59] ^ codeword[60] ^ codeword[61] ^ codeword[62] ^ codeword[63] ^ codeword[64] ^ codeword[65] ^ codeword[66] ^ codeword[67] ^ codeword[68] ^ codeword[69] ^ codeword[70] ^ codeword[71] ^ codeword[72] ^ codeword[73] ^ codeword[74] ^ codeword[75] ^ codeword[76] ^ codeword[77] ^ codeword[78] ^ codeword[79] ^ codeword[80] ^ codeword[81] ^ codeword[82] ^ codeword[83] ^ codeword[112] ^ codeword[113] ^ codeword[114] ^ codeword[115] ^ codeword[116] ^ codeword[117] ^ codeword[118] ^ codeword[119] ^ codeword[176] ^ codeword[177] ^ codeword[178] ^ codeword[179] ^ codeword[180] ^ codeword[181] ^ codeword[182] ^ codeword[183] ^ codeword[184] ^ codeword[185] ^ codeword[186] ^ codeword[187] ^ codeword[188] ^ codeword[189] ^ codeword[190] ^ codeword[191] ^ codeword[192] ^ codeword[193] ^ codeword[194] ^ codeword[195] ^ codeword[196] ^ codeword[197] ^ codeword[198] ^ codeword[199] ^ codeword[200] ^ codeword[201] ^ codeword[202] ^ codeword[203] ^ codeword[204] ^ codeword[205] ^ codeword[206] ^ codeword[207] ^ codeword[208] ^ codeword[209] ^ codeword[210] ^ codeword[211] ^ codeword[212] ^ codeword[213] ^ codeword[214] ^ codeword[215] ^ codeword[216] ^ codeword[217] ^ codeword[218] ^ codeword[219] ^ codeword[220] ^ codeword[221] ^ codeword[222] ^ codeword[223] ^ codeword[224] ^ codeword[225] ^ codeword[226] ^ codeword[227] ^ codeword[228] ^ codeword[229] ^ codeword[230] ^ codeword[231] ^ codeword[232] ^ codeword[233] ^ codeword[234] ^ codeword[235] ^ codeword[236] ^ codeword[237] ^ codeword[238] ^ codeword[239] ^ codeword[240] ^ codeword[241] ^ codeword[242] ^ codeword[243] ^ codeword[244] ^ codeword[245] ^ codeword[257];
    assign syndrome[2] = codeword[35] ^ codeword[36] ^ codeword[37] ^ codeword[38] ^ codeword[39] ^ codeword[40] ^ codeword[41] ^ codeword[42] ^ codeword[43] ^ codeword[44] ^ codeword[45] ^ codeword[46] ^ codeword[47] ^ codeword[48] ^ codeword[49] ^ codeword[50] ^ codeword[51] ^ codeword[52] ^ codeword[53] ^ codeword[54] ^ codeword[55] ^ codeword[77] ^ codeword[78] ^ codeword[79] ^ codeword[80] ^ codeword[81] ^ codeword[82] ^ codeword[83] ^ codeword[105] ^ codeword[106] ^ codeword[107] ^ codeword[108] ^ codeword[109] ^ codeword[110] ^ codeword[111] ^ codeword[119] ^ codeword[141] ^ codeword[142] ^ codeword[143] ^ codeword[144] ^ codeword[145] ^ codeword[146] ^ codeword[147] ^ codeword[148] ^ codeword[149] ^ codeword[150] ^ codeword[151] ^ codeword[152] ^ codeword[153] ^ codeword[154] ^ codeword[155] ^ codeword[156] ^ codeword[157] ^ codeword[158] ^ codeword[159] ^ codeword[160] ^ codeword[161] ^ codeword[162] ^ codeword[163] ^ codeword[164] ^ codeword[165] ^ codeword[166] ^ codeword[167] ^ codeword[168] ^ codeword[169] ^ codeword[170] ^ codeword[171] ^ codeword[172] ^ codeword[173] ^ codeword[174] ^ codeword[175] ^ codeword[211] ^ codeword[212] ^ codeword[213] ^ codeword[214] ^ codeword[215] ^ codeword[216] ^ codeword[217] ^ codeword[218] ^ codeword[219] ^ codeword[220] ^ codeword[221] ^ codeword[222] ^ codeword[223] ^ codeword[224] ^ codeword[225] ^ codeword[226] ^ codeword[227] ^ codeword[228] ^ codeword[229] ^ codeword[230] ^ codeword[231] ^ codeword[232] ^ codeword[233] ^ codeword[234] ^ codeword[235] ^ codeword[236] ^ codeword[237] ^ codeword[238] ^ codeword[239] ^ codeword[240] ^ codeword[241] ^ codeword[242] ^ codeword[243] ^ codeword[244] ^ codeword[245] ^ codeword[258];
    assign syndrome[3] = codeword[20] ^ codeword[21] ^ codeword[22] ^ codeword[23] ^ codeword[24] ^ codeword[25] ^ codeword[26] ^ codeword[27] ^ codeword[28] ^ codeword[29] ^ codeword[30] ^ codeword[31] ^ codeword[32] ^ codeword[33] ^ codeword[34] ^ codeword[50] ^ codeword[51] ^ codeword[52] ^ codeword[53] ^ codeword[54] ^ codeword[55] ^ codeword[71] ^ codeword[72] ^ codeword[73] ^ codeword[74] ^ codeword[75] ^ codeword[76] ^ codeword[83] ^ codeword[99] ^ codeword[100] ^ codeword[101] ^ codeword[102] ^ codeword[103] ^ codeword[104] ^ codeword[111] ^ codeword[118] ^ codeword[126] ^ codeword[127] ^ codeword[128] ^ codeword[129] ^ codeword[130] ^ codeword[131] ^ codeword[132] ^ codeword[133] ^ codeword[134] ^ codeword[135] ^ codeword[136] ^ codeword[137] ^ codeword[138] ^ codeword[139] ^ codeword[140] ^ codeword[156] ^ codeword[157] ^ codeword[158] ^ codeword[159] ^ codeword[160] ^ codeword[161] ^ codeword[162] ^ codeword[163] ^ codeword[164] ^ codeword[165] ^ codeword[166] ^ codeword[167] ^ codeword[168] ^ codeword[169] ^ codeword[170] ^ codeword[171] ^ codeword[172] ^ codeword[173] ^ codeword[174] ^ codeword[175] ^ codeword[191] ^ codeword[192] ^ codeword[193] ^ codeword[194] ^ codeword[195] ^ codeword[196] ^ codeword[197] ^ codeword[198] ^ codeword[199] ^ codeword[200] ^ codeword[201] ^ codeword[202] ^ codeword[203] ^ codeword[204] ^ codeword[205] ^ codeword[206] ^ codeword[207] ^ codeword[208] ^ codeword[209] ^ codeword[210] ^ codeword[231] ^ codeword[232] ^ codeword[233] ^ codeword[234] ^ codeword[235] ^ codeword[236] ^ codeword[237] ^ codeword[238] ^ codeword[239] ^ codeword[240] ^ codeword[241] ^ codeword[242] ^ codeword[243] ^ codeword[244] ^ codeword[245] ^ codeword[259];
    assign syndrome[4] = codeword[10] ^ codeword[11] ^ codeword[12] ^ codeword[13] ^ codeword[14] ^ codeword[15] ^ codeword[16] ^ codeword[17] ^ codeword[18] ^ codeword[19] ^ codeword[30] ^ codeword[31] ^ codeword[32] ^ codeword[33] ^ codeword[34] ^ codeword[45] ^ codeword[46] ^ codeword[47] ^ codeword[48] ^ codeword[49] ^ codeword[55] ^ codeword[66] ^ codeword[67] ^ codeword[68] ^ codeword[69] ^ codeword[70] ^ codeword[76] ^ codeword[82] ^ codeword[94] ^ codeword[95] ^ codeword[96] ^ codeword[97] ^ codeword[98] ^ codeword[104] ^ codeword[110] ^ codeword[117] ^ codeword[121] ^ codeword[122] ^ codeword[123] ^ codeword[124] ^ codeword[125] ^ codeword[131] ^ codeword[132] ^ codeword[133] ^ codeword[134] ^ codeword[135] ^ codeword[136] ^ codeword[137] ^ codeword[138] ^ codeword[139] ^ codeword[140] ^ codeword[146] ^ codeword[147] ^ codeword[148] ^ codeword[149] ^ codeword[150] ^ codeword[151] ^ codeword[152] ^ codeword[153] ^ codeword[154] ^ codeword[155] ^ codeword[166] ^ codeword[167] ^ codeword[168] ^ codeword[169] ^ codeword[170] ^ codeword[171] ^ codeword[172] ^ codeword[173] ^ codeword[174] ^ codeword[175] ^ codeword[181] ^ codeword[182] ^ codeword[183] ^ codeword[184] ^ codeword[185] ^ codeword[186] ^ codeword[187] ^ codeword[188] ^ codeword[189] ^ codeword[190] ^ codeword[201] ^ codeword[202] ^ codeword[203] ^ codeword[204] ^ codeword[205] ^ codeword[206] ^ codeword[207] ^ codeword[208] ^ codeword[209] ^ codeword[210] ^ codeword[221] ^ codeword[222] ^ codeword[223] ^ codeword[224] ^ codeword[225] ^ codeword[226] ^ codeword[227] ^ codeword[228] ^ codeword[229] ^ codeword[230] ^ codeword[241] ^ codeword[242] ^ codeword[243] ^ codeword[244] ^ codeword[245] ^ codeword[251] ^ codeword[252] ^ codeword[253] ^ codeword[254] ^ codeword[255] ^ codeword[260];
    assign syndrome[5] = codeword[4] ^ codeword[5] ^ codeword[6] ^ codeword[7] ^ codeword[8] ^ codeword[9] ^ codeword[16] ^ codeword[17] ^ codeword[18] ^ codeword[19] ^ codeword[26] ^ codeword[27] ^ codeword[28] ^ codeword[29] ^ codeword[34] ^ codeword[41] ^ codeword[42] ^ codeword[43] ^ codeword[44] ^ codeword[49] ^ codeword[54] ^ codeword[62] ^ codeword[63] ^ codeword[64] ^ codeword[65] ^ codeword[70] ^ codeword[75] ^ codeword[81] ^ codeword[90] ^ codeword[91] ^ codeword[92] ^ codeword[93] ^ codeword[98] ^ codeword[103] ^ codeword[109] ^ codeword[116] ^ codeword[120] ^ codeword[122] ^ codeword[123] ^ codeword[124] ^ codeword[125] ^ codeword[127] ^ codeword[128] ^ codeword[129] ^ codeword[130] ^ codeword[135] ^ codeword[136] ^ codeword[137] ^ codeword[138] ^ codeword[139] ^ codeword[140] ^ codeword[142] ^ codeword[143] ^ codeword[144] ^ codeword[145] ^ codeword[150] ^ codeword[151] ^ codeword[152] ^ codeword[153] ^ codeword[154] ^ codeword[155] ^ codeword[160] ^ codeword[161] ^ codeword[162] ^ codeword[163] ^ codeword[164] ^ codeword[165] ^ codeword[172] ^ codeword[173] ^ codeword[174] ^ codeword[175] ^ codeword[177] ^ codeword[178] ^ codeword[179] ^ codeword[180] ^ codeword[185] ^ codeword[186] ^ codeword[187] ^ codeword[188] ^ codeword[189] ^ codeword[190] ^ codeword[195] ^ codeword[196] ^ codeword[197] ^ codeword[198] ^ codeword[199] ^ codeword[200] ^ codeword[207] ^ codeword[208] ^ codeword[209] ^ codeword[210] ^ codeword[215] ^ codeword[216] ^ codeword[217] ^ codeword[218] ^ codeword[219] ^ codeword[220] ^ codeword[227] ^ codeword[228] ^ codeword[229] ^ codeword[230] ^ codeword[237] ^ codeword[238] ^ codeword[239] ^ codeword[240] ^ codeword[245] ^ codeword[247] ^ codeword[248] ^ codeword[249] ^ codeword[250] ^ codeword[255] ^ codeword[261];
    assign syndrome[6] = codeword[1] ^ codeword[2] ^ codeword[3] ^ codeword[7] ^ codeword[8] ^ codeword[9] ^ codeword[13] ^ codeword[14] ^ codeword[15] ^ codeword[19] ^ codeword[23] ^ codeword[24] ^ codeword[25] ^ codeword[29] ^ codeword[33] ^ codeword[38] ^ codeword[39] ^ codeword[40] ^ codeword[44] ^ codeword[48] ^ codeword[53] ^ codeword[59] ^ codeword[60] ^ codeword[61] ^ codeword[65] ^ codeword[69] ^ codeword[74] ^ codeword[80] ^ codeword[87] ^ codeword[88] ^ codeword[89] ^ codeword[93] ^ codeword[97] ^ codeword[102] ^ codeword[108] ^ codeword[115] ^ codeword[120] ^ codeword[121] ^ codeword[123] ^ codeword[124] ^ codeword[125] ^ codeword[126] ^ codeword[128] ^ codeword[129] ^ codeword[130] ^ codeword[132] ^ codeword[133] ^ codeword[134] ^ codeword[138] ^ codeword[139] ^ codeword[140] ^ codeword[141] ^ codeword[143] ^ codeword[144] ^ codeword[145] ^ codeword[147] ^ codeword[148] ^ codeword[149] ^ codeword[153] ^ codeword[154] ^ codeword[155] ^ codeword[157] ^ codeword[158] ^ codeword[159] ^ codeword[163] ^ codeword[164] ^ codeword[165] ^ codeword[169] ^ codeword[170] ^ codeword[171] ^ codeword[175] ^ codeword[176] ^ codeword[178] ^ codeword[179] ^ codeword[180] ^ codeword[182] ^ codeword[183] ^ codeword[184] ^ codeword[188] ^ codeword[189] ^ codeword[190] ^ codeword[192] ^ codeword[193] ^ codeword[194] ^ codeword[198] ^ codeword[199] ^ codeword[200] ^ codeword[204] ^ codeword[205] ^ codeword[206] ^ codeword[210] ^ codeword[212] ^ codeword[213] ^ codeword[214] ^ codeword[218] ^ codeword[219] ^ codeword[220] ^ codeword[224] ^ codeword[225] ^ codeword[226] ^ codeword[230] ^ codeword[234] ^ codeword[235] ^ codeword[236] ^ codeword[240] ^ codeword[244] ^ codeword[246] ^ codeword[248] ^ codeword[249] ^ codeword[250] ^ codeword[252] ^ codeword[253] ^ codeword[254] ^ codeword[262];
    assign syndrome[7] = codeword[0] ^ codeword[2] ^ codeword[3] ^ codeword[5] ^ codeword[6] ^ codeword[9] ^ codeword[11] ^ codeword[12] ^ codeword[15] ^ codeword[18] ^ codeword[21] ^ codeword[22] ^ codeword[25] ^ codeword[28] ^ codeword[32] ^ codeword[36] ^ codeword[37] ^ codeword[40] ^ codeword[43] ^ codeword[47] ^ codeword[52] ^ codeword[57] ^ codeword[58] ^ codeword[61] ^ codeword[64] ^ codeword[68] ^ codeword[73] ^ codeword[79] ^ codeword[85] ^ codeword[86] ^ codeword[89] ^ codeword[92] ^ codeword[96] ^ codeword[101] ^ codeword[107] ^ codeword[114] ^ codeword[120] ^ codeword[121] ^ codeword[122] ^ codeword[124] ^ codeword[125] ^ codeword[126] ^ codeword[127] ^ codeword[129] ^ codeword[130] ^ codeword[131] ^ codeword[133] ^ codeword[134] ^ codeword[136] ^ codeword[137] ^ codeword[140] ^ codeword[141] ^ codeword[142] ^ codeword[144] ^ codeword[145] ^ codeword[146] ^ codeword[148] ^ codeword[149] ^ codeword[151] ^ codeword[152] ^ codeword[155] ^ codeword[156] ^ codeword[158] ^ codeword[159] ^ codeword[161] ^ codeword[162] ^ codeword[165] ^ codeword[167] ^ codeword[168] ^ codeword[171] ^ codeword[174] ^ codeword[176] ^ codeword[177] ^ codeword[179] ^ codeword[180] ^ codeword[181] ^ codeword[183] ^ codeword[184] ^ codeword[186] ^ codeword[187] ^ codeword[190] ^ codeword[191] ^ codeword[193] ^ codeword[194] ^ codeword[196] ^ codeword[197] ^ codeword[200] ^ codeword[202] ^ codeword[203] ^ codeword[206] ^ codeword[209] ^ codeword[211] ^ codeword[213] ^ codeword[214] ^ codeword[216] ^ codeword[217] ^ codeword[220] ^ codeword[222] ^ codeword[223] ^ codeword[226] ^ codeword[229] ^ codeword[232] ^ codeword[233] ^ codeword[236] ^ codeword[239] ^ codeword[243] ^ codeword[246] ^ codeword[247] ^ codeword[249] ^ codeword[250] ^ codeword[251] ^ codeword[253] ^ codeword[254] ^ codeword[263];
    assign syndrome[8] = codeword[0] ^ codeword[1] ^ codeword[3] ^ codeword[4] ^ codeword[6] ^ codeword[8] ^ codeword[10] ^ codeword[12] ^ codeword[14] ^ codeword[17] ^ codeword[20] ^ codeword[22] ^ codeword[24] ^ codeword[27] ^ codeword[31] ^ codeword[35] ^ codeword[37] ^ codeword[39] ^ codeword[42] ^ codeword[46] ^ codeword[51] ^ codeword[56] ^ codeword[58] ^ codeword[60] ^ codeword[63] ^ codeword[67] ^ codeword[72] ^ codeword[78] ^ codeword[84] ^ codeword[86] ^ codeword[88] ^ codeword[91] ^ codeword[95] ^ codeword[100] ^ codeword[106] ^ codeword[113] ^ codeword[120] ^ codeword[121] ^ codeword[122] ^ codeword[123] ^ codeword[125] ^ codeword[126] ^ codeword[127] ^ codeword[128] ^ codeword[130] ^ codeword[131] ^ codeword[132] ^ codeword[134] ^ codeword[135] ^ codeword[137] ^ codeword[139] ^ codeword[141] ^ codeword[142] ^ codeword[143] ^ codeword[145] ^ codeword[146] ^ codeword[147] ^ codeword[149] ^ codeword[150] ^ codeword[152] ^ codeword[154] ^ codeword[156] ^ codeword[157] ^ codeword[159] ^ codeword[160] ^ codeword[162] ^ codeword[164] ^ codeword[166] ^ codeword[168] ^ codeword[170] ^ codeword[173] ^ codeword[176] ^ codeword[177] ^ codeword[178] ^ codeword[180] ^ codeword[181] ^ codeword[182] ^ codeword[184] ^ codeword[185] ^ codeword[187] ^ codeword[189] ^ codeword[191] ^ codeword[192] ^ codeword[194] ^ codeword[195] ^ codeword[197] ^ codeword[199] ^ codeword[201] ^ codeword[203] ^ codeword[205] ^ codeword[208] ^ codeword[211] ^ codeword[212] ^ codeword[214] ^ codeword[215] ^ codeword[217] ^ codeword[219] ^ codeword[221] ^ codeword[223] ^ codeword[225] ^ codeword[228] ^ codeword[231] ^ codeword[233] ^ codeword[235] ^ codeword[238] ^ codeword[242] ^ codeword[246] ^ codeword[247] ^ codeword[248] ^ codeword[250] ^ codeword[251] ^ codeword[252] ^ codeword[254] ^ codeword[255] ^ codeword[264];
    assign syndrome[9] = codeword[0] ^ codeword[1] ^ codeword[2] ^ codeword[4] ^ codeword[5] ^ codeword[7] ^ codeword[10] ^ codeword[11] ^ codeword[13] ^ codeword[16] ^ codeword[20] ^ codeword[21] ^ codeword[23] ^ codeword[26] ^ codeword[30] ^ codeword[35] ^ codeword[36] ^ codeword[38] ^ codeword[41] ^ codeword[45] ^ codeword[50] ^ codeword[56] ^ codeword[57] ^ codeword[59] ^ codeword[62] ^ codeword[66] ^ codeword[71] ^ codeword[77] ^ codeword[84] ^ codeword[85] ^ codeword[87] ^ codeword[90] ^ codeword[94] ^ codeword[99] ^ codeword[105] ^ codeword[112] ^ codeword[120] ^ codeword[121] ^ codeword[122] ^ codeword[123] ^ codeword[124] ^ codeword[126] ^ codeword[127] ^ codeword[128] ^ codeword[129] ^ codeword[131] ^ codeword[132] ^ codeword[133] ^ codeword[135] ^ codeword[136] ^ codeword[138] ^ codeword[141] ^ codeword[142] ^ codeword[143] ^ codeword[144] ^ codeword[146] ^ codeword[147] ^ codeword[148] ^ codeword[150] ^ codeword[151] ^ codeword[153] ^ codeword[156] ^ codeword[157] ^ codeword[158] ^ codeword[160] ^ codeword[161] ^ codeword[163] ^ codeword[166] ^ codeword[167] ^ codeword[169] ^ codeword[172] ^ codeword[176] ^ codeword[177] ^ codeword[178] ^ codeword[179] ^ codeword[181] ^ codeword[182] ^ codeword[183] ^ codeword[185] ^ codeword[186] ^ codeword[188] ^ codeword[191] ^ codeword[192] ^ codeword[193] ^ codeword[195] ^ codeword[196] ^ codeword[198] ^ codeword[201] ^ codeword[202] ^ codeword[204] ^ codeword[207] ^ codeword[211] ^ codeword[212] ^ codeword[213] ^ codeword[215] ^ codeword[216] ^ codeword[218] ^ codeword[221] ^ codeword[222] ^ codeword[224] ^ codeword[227] ^ codeword[231] ^ codeword[232] ^ codeword[234] ^ codeword[237] ^ codeword[241] ^ codeword[246] ^ codeword[247] ^ codeword[248] ^ codeword[249] ^ codeword[251] ^ codeword[252] ^ codeword[253] ^ codeword[255] ^ codeword[265];
  end else if (CodewordWidth == 523 && MessageWidth == 512) begin : gen_523_512
    `BR_ASSERT_STATIC(parity_width_matches_a, ParityWidth == 11)
    assign syndrome[0] = codeword[120] ^ codeword[121] ^ codeword[122] ^ codeword[123] ^ codeword[124] ^ codeword[125] ^ codeword[126] ^ codeword[127] ^ codeword[128] ^ codeword[129] ^ codeword[130] ^ codeword[131] ^ codeword[132] ^ codeword[133] ^ codeword[134] ^ codeword[135] ^ codeword[136] ^ codeword[137] ^ codeword[138] ^ codeword[139] ^ codeword[140] ^ codeword[141] ^ codeword[142] ^ codeword[143] ^ codeword[144] ^ codeword[145] ^ codeword[146] ^ codeword[147] ^ codeword[148] ^ codeword[149] ^ codeword[150] ^ codeword[151] ^ codeword[152] ^ codeword[153] ^ codeword[154] ^ codeword[155] ^ codeword[156] ^ codeword[157] ^ codeword[158] ^ codeword[159] ^ codeword[160] ^ codeword[161] ^ codeword[162] ^ codeword[163] ^ codeword[164] ^ codeword[417] ^ codeword[418] ^ codeword[419] ^ codeword[420] ^ codeword[421] ^ codeword[422] ^ codeword[423] ^ codeword[424] ^ codeword[425] ^ codeword[426] ^ codeword[427] ^ codeword[428] ^ codeword[429] ^ codeword[430] ^ codeword[431] ^ codeword[432] ^ codeword[433] ^ codeword[434] ^ codeword[435] ^ codeword[436] ^ codeword[437] ^ codeword[438] ^ codeword[439] ^ codeword[440] ^ codeword[441] ^ codeword[442] ^ codeword[443] ^ codeword[444] ^ codeword[445] ^ codeword[446] ^ codeword[447] ^ codeword[448] ^ codeword[449] ^ codeword[450] ^ codeword[451] ^ codeword[452] ^ codeword[453] ^ codeword[454] ^ codeword[455] ^ codeword[456] ^ codeword[457] ^ codeword[458] ^ codeword[459] ^ codeword[460] ^ codeword[461] ^ codeword[462] ^ codeword[463] ^ codeword[464] ^ codeword[465] ^ codeword[466] ^ codeword[467] ^ codeword[468] ^ codeword[469] ^ codeword[470] ^ codeword[471] ^ codeword[472] ^ codeword[473] ^ codeword[474] ^ codeword[475] ^ codeword[476] ^ codeword[477] ^ codeword[478] ^ codeword[479] ^ codeword[480] ^ codeword[481] ^ codeword[482] ^ codeword[483] ^ codeword[484] ^ codeword[485] ^ codeword[486] ^ codeword[487] ^ codeword[488] ^ codeword[489] ^ codeword[490] ^ codeword[491] ^ codeword[492] ^ codeword[493] ^ codeword[494] ^ codeword[495] ^ codeword[496] ^ codeword[497] ^ codeword[498] ^ codeword[499] ^ codeword[500] ^ codeword[501] ^ codeword[502] ^ codeword[503] ^ codeword[504] ^ codeword[505] ^ codeword[506] ^ codeword[507] ^ codeword[508] ^ codeword[509] ^ codeword[510] ^ codeword[511] ^ codeword[512];
    assign syndrome[1] = codeword[84] ^ codeword[85] ^ codeword[86] ^ codeword[87] ^ codeword[88] ^ codeword[89] ^ codeword[90] ^ codeword[91] ^ codeword[92] ^ codeword[93] ^ codeword[94] ^ codeword[95] ^ codeword[96] ^ codeword[97] ^ codeword[98] ^ codeword[99] ^ codeword[100] ^ codeword[101] ^ codeword[102] ^ codeword[103] ^ codeword[104] ^ codeword[105] ^ codeword[106] ^ codeword[107] ^ codeword[108] ^ codeword[109] ^ codeword[110] ^ codeword[111] ^ codeword[112] ^ codeword[113] ^ codeword[114] ^ codeword[115] ^ codeword[116] ^ codeword[117] ^ codeword[118] ^ codeword[119] ^ codeword[156] ^ codeword[157] ^ codeword[158] ^ codeword[159] ^ codeword[160] ^ codeword[161] ^ codeword[162] ^ codeword[163] ^ codeword[164] ^ codeword[291] ^ codeword[292] ^ codeword[293] ^ codeword[294] ^ codeword[295] ^ codeword[296] ^ codeword[297] ^ codeword[298] ^ codeword[299] ^ codeword[300] ^ codeword[301] ^ codeword[302] ^ codeword[303] ^ codeword[304] ^ codeword[305] ^ codeword[306] ^ codeword[307] ^ codeword[308] ^ codeword[309] ^ codeword[310] ^ codeword[311] ^ codeword[312] ^ codeword[313] ^ codeword[314] ^ codeword[315] ^ codeword[316] ^ codeword[317] ^ codeword[318] ^ codeword[319] ^ codeword[320] ^ codeword[321] ^ codeword[322] ^ codeword[323] ^ codeword[324] ^ codeword[325] ^ codeword[326] ^ codeword[327] ^ codeword[328] ^ codeword[329] ^ codeword[330] ^ codeword[331] ^ codeword[332] ^ codeword[333] ^ codeword[334] ^ codeword[335] ^ codeword[336] ^ codeword[337] ^ codeword[338] ^ codeword[339] ^ codeword[340] ^ codeword[341] ^ codeword[342] ^ codeword[343] ^ codeword[344] ^ codeword[345] ^ codeword[346] ^ codeword[347] ^ codeword[348] ^ codeword[349] ^ codeword[350] ^ codeword[351] ^ codeword[352] ^ codeword[353] ^ codeword[354] ^ codeword[355] ^ codeword[356] ^ codeword[357] ^ codeword[358] ^ codeword[359] ^ codeword[360] ^ codeword[361] ^ codeword[362] ^ codeword[363] ^ codeword[364] ^ codeword[365] ^ codeword[366] ^ codeword[367] ^ codeword[368] ^ codeword[369] ^ codeword[370] ^ codeword[371] ^ codeword[372] ^ codeword[373] ^ codeword[374] ^ codeword[375] ^ codeword[376] ^ codeword[377] ^ codeword[378] ^ codeword[379] ^ codeword[380] ^ codeword[381] ^ codeword[382] ^ codeword[383] ^ codeword[384] ^ codeword[385] ^ codeword[386] ^ codeword[387] ^ codeword[388] ^ codeword[389] ^ codeword[390] ^ codeword[391] ^ codeword[392] ^ codeword[393] ^ codeword[394] ^ codeword[395] ^ codeword[396] ^ codeword[397] ^ codeword[398] ^ codeword[399] ^ codeword[400] ^ codeword[401] ^ codeword[402] ^ codeword[403] ^ codeword[404] ^ codeword[405] ^ codeword[406] ^ codeword[407] ^ codeword[408] ^ codeword[409] ^ codeword[410] ^ codeword[411] ^ codeword[412] ^ codeword[413] ^ codeword[414] ^ codeword[415] ^ codeword[416] ^ codeword[513];
    assign syndrome[2] = codeword[56] ^ codeword[57] ^ codeword[58] ^ codeword[59] ^ codeword[60] ^ codeword[61] ^ codeword[62] ^ codeword[63] ^ codeword[64] ^ codeword[65] ^ codeword[66] ^ codeword[67] ^ codeword[68] ^ codeword[69] ^ codeword[70] ^ codeword[71] ^ codeword[72] ^ codeword[73] ^ codeword[74] ^ codeword[75] ^ codeword[76] ^ codeword[77] ^ codeword[78] ^ codeword[79] ^ codeword[80] ^ codeword[81] ^ codeword[82] ^ codeword[83] ^ codeword[112] ^ codeword[113] ^ codeword[114] ^ codeword[115] ^ codeword[116] ^ codeword[117] ^ codeword[118] ^ codeword[119] ^ codeword[148] ^ codeword[149] ^ codeword[150] ^ codeword[151] ^ codeword[152] ^ codeword[153] ^ codeword[154] ^ codeword[155] ^ codeword[164] ^ codeword[221] ^ codeword[222] ^ codeword[223] ^ codeword[224] ^ codeword[225] ^ codeword[226] ^ codeword[227] ^ codeword[228] ^ codeword[229] ^ codeword[230] ^ codeword[231] ^ codeword[232] ^ codeword[233] ^ codeword[234] ^ codeword[235] ^ codeword[236] ^ codeword[237] ^ codeword[238] ^ codeword[239] ^ codeword[240] ^ codeword[241] ^ codeword[242] ^ codeword[243] ^ codeword[244] ^ codeword[245] ^ codeword[246] ^ codeword[247] ^ codeword[248] ^ codeword[249] ^ codeword[250] ^ codeword[251] ^ codeword[252] ^ codeword[253] ^ codeword[254] ^ codeword[255] ^ codeword[256] ^ codeword[257] ^ codeword[258] ^ codeword[259] ^ codeword[260] ^ codeword[261] ^ codeword[262] ^ codeword[263] ^ codeword[264] ^ codeword[265] ^ codeword[266] ^ codeword[267] ^ codeword[268] ^ codeword[269] ^ codeword[270] ^ codeword[271] ^ codeword[272] ^ codeword[273] ^ codeword[274] ^ codeword[275] ^ codeword[276] ^ codeword[277] ^ codeword[278] ^ codeword[279] ^ codeword[280] ^ codeword[281] ^ codeword[282] ^ codeword[283] ^ codeword[284] ^ codeword[285] ^ codeword[286] ^ codeword[287] ^ codeword[288] ^ codeword[289] ^ codeword[290] ^ codeword[361] ^ codeword[362] ^ codeword[363] ^ codeword[364] ^ codeword[365] ^ codeword[366] ^ codeword[367] ^ codeword[368] ^ codeword[369] ^ codeword[370] ^ codeword[371] ^ codeword[372] ^ codeword[373] ^ codeword[374] ^ codeword[375] ^ codeword[376] ^ codeword[377] ^ codeword[378] ^ codeword[379] ^ codeword[380] ^ codeword[381] ^ codeword[382] ^ codeword[383] ^ codeword[384] ^ codeword[385] ^ codeword[386] ^ codeword[387] ^ codeword[388] ^ codeword[389] ^ codeword[390] ^ codeword[391] ^ codeword[392] ^ codeword[393] ^ codeword[394] ^ codeword[395] ^ codeword[396] ^ codeword[397] ^ codeword[398] ^ codeword[399] ^ codeword[400] ^ codeword[401] ^ codeword[402] ^ codeword[403] ^ codeword[404] ^ codeword[405] ^ codeword[406] ^ codeword[407] ^ codeword[408] ^ codeword[409] ^ codeword[410] ^ codeword[411] ^ codeword[412] ^ codeword[413] ^ codeword[414] ^ codeword[415] ^ codeword[416] ^ codeword[487] ^ codeword[488] ^ codeword[489] ^ codeword[490] ^ codeword[491] ^ codeword[492] ^ codeword[493] ^ codeword[494] ^ codeword[495] ^ codeword[496] ^ codeword[497] ^ codeword[498] ^ codeword[499] ^ codeword[500] ^ codeword[501] ^ codeword[502] ^ codeword[503] ^ codeword[504] ^ codeword[505] ^ codeword[506] ^ codeword[507] ^ codeword[508] ^ codeword[509] ^ codeword[510] ^ codeword[511] ^ codeword[514];
    assign syndrome[3] = codeword[35] ^ codeword[36] ^ codeword[37] ^ codeword[38] ^ codeword[39] ^ codeword[40] ^ codeword[41] ^ codeword[42] ^ codeword[43] ^ codeword[44] ^ codeword[45] ^ codeword[46] ^ codeword[47] ^ codeword[48] ^ codeword[49] ^ codeword[50] ^ codeword[51] ^ codeword[52] ^ codeword[53] ^ codeword[54] ^ codeword[55] ^ codeword[77] ^ codeword[78] ^ codeword[79] ^ codeword[80] ^ codeword[81] ^ codeword[82] ^ codeword[83] ^ codeword[105] ^ codeword[106] ^ codeword[107] ^ codeword[108] ^ codeword[109] ^ codeword[110] ^ codeword[111] ^ codeword[119] ^ codeword[141] ^ codeword[142] ^ codeword[143] ^ codeword[144] ^ codeword[145] ^ codeword[146] ^ codeword[147] ^ codeword[155] ^ codeword[163] ^ codeword[186] ^ codeword[187] ^ codeword[188] ^ codeword[189] ^ codeword[190] ^ codeword[191] ^ codeword[192] ^ codeword[193] ^ codeword[194] ^ codeword[195] ^ codeword[196] ^ codeword[197] ^ codeword[198] ^ codeword[199] ^ codeword[200] ^ codeword[201] ^ codeword[202] ^ codeword[203] ^ codeword[204] ^ codeword[205] ^ codeword[206] ^ codeword[207] ^ codeword[208] ^ codeword[209] ^ codeword[210] ^ codeword[211] ^ codeword[212] ^ codeword[213] ^ codeword[214] ^ codeword[215] ^ codeword[216] ^ codeword[217] ^ codeword[218] ^ codeword[219] ^ codeword[220] ^ codeword[256] ^ codeword[257] ^ codeword[258] ^ codeword[259] ^ codeword[260] ^ codeword[261] ^ codeword[262] ^ codeword[263] ^ codeword[264] ^ codeword[265] ^ codeword[266] ^ codeword[267] ^ codeword[268] ^ codeword[269] ^ codeword[270] ^ codeword[271] ^ codeword[272] ^ codeword[273] ^ codeword[274] ^ codeword[275] ^ codeword[276] ^ codeword[277] ^ codeword[278] ^ codeword[279] ^ codeword[280] ^ codeword[281] ^ codeword[282] ^ codeword[283] ^ codeword[284] ^ codeword[285] ^ codeword[286] ^ codeword[287] ^ codeword[288] ^ codeword[289] ^ codeword[290] ^ codeword[326] ^ codeword[327] ^ codeword[328] ^ codeword[329] ^ codeword[330] ^ codeword[331] ^ codeword[332] ^ codeword[333] ^ codeword[334] ^ codeword[335] ^ codeword[336] ^ codeword[337] ^ codeword[338] ^ codeword[339] ^ codeword[340] ^ codeword[341] ^ codeword[342] ^ codeword[343] ^ codeword[344] ^ codeword[345] ^ codeword[346] ^ codeword[347] ^ codeword[348] ^ codeword[349] ^ codeword[350] ^ codeword[351] ^ codeword[352] ^ codeword[353] ^ codeword[354] ^ codeword[355] ^ codeword[356] ^ codeword[357] ^ codeword[358] ^ codeword[359] ^ codeword[360] ^ codeword[396] ^ codeword[397] ^ codeword[398] ^ codeword[399] ^ codeword[400] ^ codeword[401] ^ codeword[402] ^ codeword[403] ^ codeword[404] ^ codeword[405] ^ codeword[406] ^ codeword[407] ^ codeword[408] ^ codeword[409] ^ codeword[410] ^ codeword[411] ^ codeword[412] ^ codeword[413] ^ codeword[414] ^ codeword[415] ^ codeword[416] ^ codeword[452] ^ codeword[453] ^ codeword[454] ^ codeword[455] ^ codeword[456] ^ codeword[457] ^ codeword[458] ^ codeword[459] ^ codeword[460] ^ codeword[461] ^ codeword[462] ^ codeword[463] ^ codeword[464] ^ codeword[465] ^ codeword[466] ^ codeword[467] ^ codeword[468] ^ codeword[469] ^ codeword[470] ^ codeword[471] ^ codeword[472] ^ codeword[473] ^ codeword[474] ^ codeword[475] ^ codeword[476] ^ codeword[477] ^ codeword[478] ^ codeword[479] ^ codeword[480] ^ codeword[481] ^ codeword[482] ^ codeword[483] ^ codeword[484] ^ codeword[485] ^ codeword[486] ^ codeword[515];
    assign syndrome[4] = codeword[20] ^ codeword[21] ^ codeword[22] ^ codeword[23] ^ codeword[24] ^ codeword[25] ^ codeword[26] ^ codeword[27] ^ codeword[28] ^ codeword[29] ^ codeword[30] ^ codeword[31] ^ codeword[32] ^ codeword[33] ^ codeword[34] ^ codeword[50] ^ codeword[51] ^ codeword[52] ^ codeword[53] ^ codeword[54] ^ codeword[55] ^ codeword[71] ^ codeword[72] ^ codeword[73] ^ codeword[74] ^ codeword[75] ^ codeword[76] ^ codeword[83] ^ codeword[99] ^ codeword[100] ^ codeword[101] ^ codeword[102] ^ codeword[103] ^ codeword[104] ^ codeword[111] ^ codeword[118] ^ codeword[135] ^ codeword[136] ^ codeword[137] ^ codeword[138] ^ codeword[139] ^ codeword[140] ^ codeword[147] ^ codeword[154] ^ codeword[162] ^ codeword[171] ^ codeword[172] ^ codeword[173] ^ codeword[174] ^ codeword[175] ^ codeword[176] ^ codeword[177] ^ codeword[178] ^ codeword[179] ^ codeword[180] ^ codeword[181] ^ codeword[182] ^ codeword[183] ^ codeword[184] ^ codeword[185] ^ codeword[201] ^ codeword[202] ^ codeword[203] ^ codeword[204] ^ codeword[205] ^ codeword[206] ^ codeword[207] ^ codeword[208] ^ codeword[209] ^ codeword[210] ^ codeword[211] ^ codeword[212] ^ codeword[213] ^ codeword[214] ^ codeword[215] ^ codeword[216] ^ codeword[217] ^ codeword[218] ^ codeword[219] ^ codeword[220] ^ codeword[236] ^ codeword[237] ^ codeword[238] ^ codeword[239] ^ codeword[240] ^ codeword[241] ^ codeword[242] ^ codeword[243] ^ codeword[244] ^ codeword[245] ^ codeword[246] ^ codeword[247] ^ codeword[248] ^ codeword[249] ^ codeword[250] ^ codeword[251] ^ codeword[252] ^ codeword[253] ^ codeword[254] ^ codeword[255] ^ codeword[276] ^ codeword[277] ^ codeword[278] ^ codeword[279] ^ codeword[280] ^ codeword[281] ^ codeword[282] ^ codeword[283] ^ codeword[284] ^ codeword[285] ^ codeword[286] ^ codeword[287] ^ codeword[288] ^ codeword[289] ^ codeword[290] ^ codeword[306] ^ codeword[307] ^ codeword[308] ^ codeword[309] ^ codeword[310] ^ codeword[311] ^ codeword[312] ^ codeword[313] ^ codeword[314] ^ codeword[315] ^ codeword[316] ^ codeword[317] ^ codeword[318] ^ codeword[319] ^ codeword[320] ^ codeword[321] ^ codeword[322] ^ codeword[323] ^ codeword[324] ^ codeword[325] ^ codeword[346] ^ codeword[347] ^ codeword[348] ^ codeword[349] ^ codeword[350] ^ codeword[351] ^ codeword[352] ^ codeword[353] ^ codeword[354] ^ codeword[355] ^ codeword[356] ^ codeword[357] ^ codeword[358] ^ codeword[359] ^ codeword[360] ^ codeword[381] ^ codeword[382] ^ codeword[383] ^ codeword[384] ^ codeword[385] ^ codeword[386] ^ codeword[387] ^ codeword[388] ^ codeword[389] ^ codeword[390] ^ codeword[391] ^ codeword[392] ^ codeword[393] ^ codeword[394] ^ codeword[395] ^ codeword[411] ^ codeword[412] ^ codeword[413] ^ codeword[414] ^ codeword[415] ^ codeword[416] ^ codeword[432] ^ codeword[433] ^ codeword[434] ^ codeword[435] ^ codeword[436] ^ codeword[437] ^ codeword[438] ^ codeword[439] ^ codeword[440] ^ codeword[441] ^ codeword[442] ^ codeword[443] ^ codeword[444] ^ codeword[445] ^ codeword[446] ^ codeword[447] ^ codeword[448] ^ codeword[449] ^ codeword[450] ^ codeword[451] ^ codeword[472] ^ codeword[473] ^ codeword[474] ^ codeword[475] ^ codeword[476] ^ codeword[477] ^ codeword[478] ^ codeword[479] ^ codeword[480] ^ codeword[481] ^ codeword[482] ^ codeword[483] ^ codeword[484] ^ codeword[485] ^ codeword[486] ^ codeword[507] ^ codeword[508] ^ codeword[509] ^ codeword[510] ^ codeword[511] ^ codeword[516];
    assign syndrome[5] = codeword[10] ^ codeword[11] ^ codeword[12] ^ codeword[13] ^ codeword[14] ^ codeword[15] ^ codeword[16] ^ codeword[17] ^ codeword[18] ^ codeword[19] ^ codeword[30] ^ codeword[31] ^ codeword[32] ^ codeword[33] ^ codeword[34] ^ codeword[45] ^ codeword[46] ^ codeword[47] ^ codeword[48] ^ codeword[49] ^ codeword[55] ^ codeword[66] ^ codeword[67] ^ codeword[68] ^ codeword[69] ^ codeword[70] ^ codeword[76] ^ codeword[82] ^ codeword[94] ^ codeword[95] ^ codeword[96] ^ codeword[97] ^ codeword[98] ^ codeword[104] ^ codeword[110] ^ codeword[117] ^ codeword[130] ^ codeword[131] ^ codeword[132] ^ codeword[133] ^ codeword[134] ^ codeword[140] ^ codeword[146] ^ codeword[153] ^ codeword[161] ^ codeword[166] ^ codeword[167] ^ codeword[168] ^ codeword[169] ^ codeword[170] ^ codeword[176] ^ codeword[177] ^ codeword[178] ^ codeword[179] ^ codeword[180] ^ codeword[181] ^ codeword[182] ^ codeword[183] ^ codeword[184] ^ codeword[185] ^ codeword[191] ^ codeword[192] ^ codeword[193] ^ codeword[194] ^ codeword[195] ^ codeword[196] ^ codeword[197] ^ codeword[198] ^ codeword[199] ^ codeword[200] ^ codeword[211] ^ codeword[212] ^ codeword[213] ^ codeword[214] ^ codeword[215] ^ codeword[216] ^ codeword[217] ^ codeword[218] ^ codeword[219] ^ codeword[220] ^ codeword[226] ^ codeword[227] ^ codeword[228] ^ codeword[229] ^ codeword[230] ^ codeword[231] ^ codeword[232] ^ codeword[233] ^ codeword[234] ^ codeword[235] ^ codeword[246] ^ codeword[247] ^ codeword[248] ^ codeword[249] ^ codeword[250] ^ codeword[251] ^ codeword[252] ^ codeword[253] ^ codeword[254] ^ codeword[255] ^ codeword[266] ^ codeword[267] ^ codeword[268] ^ codeword[269] ^ codeword[270] ^ codeword[271] ^ codeword[272] ^ codeword[273] ^ codeword[274] ^ codeword[275] ^ codeword[286] ^ codeword[287] ^ codeword[288] ^ codeword[289] ^ codeword[290] ^ codeword[296] ^ codeword[297] ^ codeword[298] ^ codeword[299] ^ codeword[300] ^ codeword[301] ^ codeword[302] ^ codeword[303] ^ codeword[304] ^ codeword[305] ^ codeword[316] ^ codeword[317] ^ codeword[318] ^ codeword[319] ^ codeword[320] ^ codeword[321] ^ codeword[322] ^ codeword[323] ^ codeword[324] ^ codeword[325] ^ codeword[336] ^ codeword[337] ^ codeword[338] ^ codeword[339] ^ codeword[340] ^ codeword[341] ^ codeword[342] ^ codeword[343] ^ codeword[344] ^ codeword[345] ^ codeword[356] ^ codeword[357] ^ codeword[358] ^ codeword[359] ^ codeword[360] ^ codeword[371] ^ codeword[372] ^ codeword[373] ^ codeword[374] ^ codeword[375] ^ codeword[376] ^ codeword[377] ^ codeword[378] ^ codeword[379] ^ codeword[380] ^ codeword[391] ^ codeword[392] ^ codeword[393] ^ codeword[394] ^ codeword[395] ^ codeword[406] ^ codeword[407] ^ codeword[408] ^ codeword[409] ^ codeword[410] ^ codeword[416] ^ codeword[422] ^ codeword[423] ^ codeword[424] ^ codeword[425] ^ codeword[426] ^ codeword[427] ^ codeword[428] ^ codeword[429] ^ codeword[430] ^ codeword[431] ^ codeword[442] ^ codeword[443] ^ codeword[444] ^ codeword[445] ^ codeword[446] ^ codeword[447] ^ codeword[448] ^ codeword[449] ^ codeword[450] ^ codeword[451] ^ codeword[462] ^ codeword[463] ^ codeword[464] ^ codeword[465] ^ codeword[466] ^ codeword[467] ^ codeword[468] ^ codeword[469] ^ codeword[470] ^ codeword[471] ^ codeword[482] ^ codeword[483] ^ codeword[484] ^ codeword[485] ^ codeword[486] ^ codeword[497] ^ codeword[498] ^ codeword[499] ^ codeword[500] ^ codeword[501] ^ codeword[502] ^ codeword[503] ^ codeword[504] ^ codeword[505] ^ codeword[506] ^ codeword[517];
    assign syndrome[6] = codeword[4] ^ codeword[5] ^ codeword[6] ^ codeword[7] ^ codeword[8] ^ codeword[9] ^ codeword[16] ^ codeword[17] ^ codeword[18] ^ codeword[19] ^ codeword[26] ^ codeword[27] ^ codeword[28] ^ codeword[29] ^ codeword[34] ^ codeword[41] ^ codeword[42] ^ codeword[43] ^ codeword[44] ^ codeword[49] ^ codeword[54] ^ codeword[62] ^ codeword[63] ^ codeword[64] ^ codeword[65] ^ codeword[70] ^ codeword[75] ^ codeword[81] ^ codeword[90] ^ codeword[91] ^ codeword[92] ^ codeword[93] ^ codeword[98] ^ codeword[103] ^ codeword[109] ^ codeword[116] ^ codeword[126] ^ codeword[127] ^ codeword[128] ^ codeword[129] ^ codeword[134] ^ codeword[139] ^ codeword[145] ^ codeword[152] ^ codeword[160] ^ codeword[165] ^ codeword[167] ^ codeword[168] ^ codeword[169] ^ codeword[170] ^ codeword[172] ^ codeword[173] ^ codeword[174] ^ codeword[175] ^ codeword[180] ^ codeword[181] ^ codeword[182] ^ codeword[183] ^ codeword[184] ^ codeword[185] ^ codeword[187] ^ codeword[188] ^ codeword[189] ^ codeword[190] ^ codeword[195] ^ codeword[196] ^ codeword[197] ^ codeword[198] ^ codeword[199] ^ codeword[200] ^ codeword[205] ^ codeword[206] ^ codeword[207] ^ codeword[208] ^ codeword[209] ^ codeword[210] ^ codeword[217] ^ codeword[218] ^ codeword[219] ^ codeword[220] ^ codeword[222] ^ codeword[223] ^ codeword[224] ^ codeword[225] ^ codeword[230] ^ codeword[231] ^ codeword[232] ^ codeword[233] ^ codeword[234] ^ codeword[235] ^ codeword[240] ^ codeword[241] ^ codeword[242] ^ codeword[243] ^ codeword[244] ^ codeword[245] ^ codeword[252] ^ codeword[253] ^ codeword[254] ^ codeword[255] ^ codeword[260] ^ codeword[261] ^ codeword[262] ^ codeword[263] ^ codeword[264] ^ codeword[265] ^ codeword[272] ^ codeword[273] ^ codeword[274] ^ codeword[275] ^ codeword[282] ^ codeword[283] ^ codeword[284] ^ codeword[285] ^ codeword[290] ^ codeword[292] ^ codeword[293] ^ codeword[294] ^ codeword[295] ^ codeword[300] ^ codeword[301] ^ codeword[302] ^ codeword[303] ^ codeword[304] ^ codeword[305] ^ codeword[310] ^ codeword[311] ^ codeword[312] ^ codeword[313] ^ codeword[314] ^ codeword[315] ^ codeword[322] ^ codeword[323] ^ codeword[324] ^ codeword[325] ^ codeword[330] ^ codeword[331] ^ codeword[332] ^ codeword[333] ^ codeword[334] ^ codeword[335] ^ codeword[342] ^ codeword[343] ^ codeword[344] ^ codeword[345] ^ codeword[352] ^ codeword[353] ^ codeword[354] ^ codeword[355] ^ codeword[360] ^ codeword[365] ^ codeword[366] ^ codeword[367] ^ codeword[368] ^ codeword[369] ^ codeword[370] ^ codeword[377] ^ codeword[378] ^ codeword[379] ^ codeword[380] ^ codeword[387] ^ codeword[388] ^ codeword[389] ^ codeword[390] ^ codeword[395] ^ codeword[402] ^ codeword[403] ^ codeword[404] ^ codeword[405] ^ codeword[410] ^ codeword[415] ^ codeword[418] ^ codeword[419] ^ codeword[420] ^ codeword[421] ^ codeword[426] ^ codeword[427] ^ codeword[428] ^ codeword[429] ^ codeword[430] ^ codeword[431] ^ codeword[436] ^ codeword[437] ^ codeword[438] ^ codeword[439] ^ codeword[440] ^ codeword[441] ^ codeword[448] ^ codeword[449] ^ codeword[450] ^ codeword[451] ^ codeword[456] ^ codeword[457] ^ codeword[458] ^ codeword[459] ^ codeword[460] ^ codeword[461] ^ codeword[468] ^ codeword[469] ^ codeword[470] ^ codeword[471] ^ codeword[478] ^ codeword[479] ^ codeword[480] ^ codeword[481] ^ codeword[486] ^ codeword[491] ^ codeword[492] ^ codeword[493] ^ codeword[494] ^ codeword[495] ^ codeword[496] ^ codeword[503] ^ codeword[504] ^ codeword[505] ^ codeword[506] ^ codeword[518];
    assign syndrome[7] = codeword[1] ^ codeword[2] ^ codeword[3] ^ codeword[7] ^ codeword[8] ^ codeword[9] ^ codeword[13] ^ codeword[14] ^ codeword[15] ^ codeword[19] ^ codeword[23] ^ codeword[24] ^ codeword[25] ^ codeword[29] ^ codeword[33] ^ codeword[38] ^ codeword[39] ^ codeword[40] ^ codeword[44] ^ codeword[48] ^ codeword[53] ^ codeword[59] ^ codeword[60] ^ codeword[61] ^ codeword[65] ^ codeword[69] ^ codeword[74] ^ codeword[80] ^ codeword[87] ^ codeword[88] ^ codeword[89] ^ codeword[93] ^ codeword[97] ^ codeword[102] ^ codeword[108] ^ codeword[115] ^ codeword[123] ^ codeword[124] ^ codeword[125] ^ codeword[129] ^ codeword[133] ^ codeword[138] ^ codeword[144] ^ codeword[151] ^ codeword[159] ^ codeword[165] ^ codeword[166] ^ codeword[168] ^ codeword[169] ^ codeword[170] ^ codeword[171] ^ codeword[173] ^ codeword[174] ^ codeword[175] ^ codeword[177] ^ codeword[178] ^ codeword[179] ^ codeword[183] ^ codeword[184] ^ codeword[185] ^ codeword[186] ^ codeword[188] ^ codeword[189] ^ codeword[190] ^ codeword[192] ^ codeword[193] ^ codeword[194] ^ codeword[198] ^ codeword[199] ^ codeword[200] ^ codeword[202] ^ codeword[203] ^ codeword[204] ^ codeword[208] ^ codeword[209] ^ codeword[210] ^ codeword[214] ^ codeword[215] ^ codeword[216] ^ codeword[220] ^ codeword[221] ^ codeword[223] ^ codeword[224] ^ codeword[225] ^ codeword[227] ^ codeword[228] ^ codeword[229] ^ codeword[233] ^ codeword[234] ^ codeword[235] ^ codeword[237] ^ codeword[238] ^ codeword[239] ^ codeword[243] ^ codeword[244] ^ codeword[245] ^ codeword[249] ^ codeword[250] ^ codeword[251] ^ codeword[255] ^ codeword[257] ^ codeword[258] ^ codeword[259] ^ codeword[263] ^ codeword[264] ^ codeword[265] ^ codeword[269] ^ codeword[270] ^ codeword[271] ^ codeword[275] ^ codeword[279] ^ codeword[280] ^ codeword[281] ^ codeword[285] ^ codeword[289] ^ codeword[291] ^ codeword[293] ^ codeword[294] ^ codeword[295] ^ codeword[297] ^ codeword[298] ^ codeword[299] ^ codeword[303] ^ codeword[304] ^ codeword[305] ^ codeword[307] ^ codeword[308] ^ codeword[309] ^ codeword[313] ^ codeword[314] ^ codeword[315] ^ codeword[319] ^ codeword[320] ^ codeword[321] ^ codeword[325] ^ codeword[327] ^ codeword[328] ^ codeword[329] ^ codeword[333] ^ codeword[334] ^ codeword[335] ^ codeword[339] ^ codeword[340] ^ codeword[341] ^ codeword[345] ^ codeword[349] ^ codeword[350] ^ codeword[351] ^ codeword[355] ^ codeword[359] ^ codeword[362] ^ codeword[363] ^ codeword[364] ^ codeword[368] ^ codeword[369] ^ codeword[370] ^ codeword[374] ^ codeword[375] ^ codeword[376] ^ codeword[380] ^ codeword[384] ^ codeword[385] ^ codeword[386] ^ codeword[390] ^ codeword[394] ^ codeword[399] ^ codeword[400] ^ codeword[401] ^ codeword[405] ^ codeword[409] ^ codeword[414] ^ codeword[417] ^ codeword[419] ^ codeword[420] ^ codeword[421] ^ codeword[423] ^ codeword[424] ^ codeword[425] ^ codeword[429] ^ codeword[430] ^ codeword[431] ^ codeword[433] ^ codeword[434] ^ codeword[435] ^ codeword[439] ^ codeword[440] ^ codeword[441] ^ codeword[445] ^ codeword[446] ^ codeword[447] ^ codeword[451] ^ codeword[453] ^ codeword[454] ^ codeword[455] ^ codeword[459] ^ codeword[460] ^ codeword[461] ^ codeword[465] ^ codeword[466] ^ codeword[467] ^ codeword[471] ^ codeword[475] ^ codeword[476] ^ codeword[477] ^ codeword[481] ^ codeword[485] ^ codeword[488] ^ codeword[489] ^ codeword[490] ^ codeword[494] ^ codeword[495] ^ codeword[496] ^ codeword[500] ^ codeword[501] ^ codeword[502] ^ codeword[506] ^ codeword[510] ^ codeword[511] ^ codeword[519];
    assign syndrome[8] = codeword[0] ^ codeword[2] ^ codeword[3] ^ codeword[5] ^ codeword[6] ^ codeword[9] ^ codeword[11] ^ codeword[12] ^ codeword[15] ^ codeword[18] ^ codeword[21] ^ codeword[22] ^ codeword[25] ^ codeword[28] ^ codeword[32] ^ codeword[36] ^ codeword[37] ^ codeword[40] ^ codeword[43] ^ codeword[47] ^ codeword[52] ^ codeword[57] ^ codeword[58] ^ codeword[61] ^ codeword[64] ^ codeword[68] ^ codeword[73] ^ codeword[79] ^ codeword[85] ^ codeword[86] ^ codeword[89] ^ codeword[92] ^ codeword[96] ^ codeword[101] ^ codeword[107] ^ codeword[114] ^ codeword[121] ^ codeword[122] ^ codeword[125] ^ codeword[128] ^ codeword[132] ^ codeword[137] ^ codeword[143] ^ codeword[150] ^ codeword[158] ^ codeword[165] ^ codeword[166] ^ codeword[167] ^ codeword[169] ^ codeword[170] ^ codeword[171] ^ codeword[172] ^ codeword[174] ^ codeword[175] ^ codeword[176] ^ codeword[178] ^ codeword[179] ^ codeword[181] ^ codeword[182] ^ codeword[185] ^ codeword[186] ^ codeword[187] ^ codeword[189] ^ codeword[190] ^ codeword[191] ^ codeword[193] ^ codeword[194] ^ codeword[196] ^ codeword[197] ^ codeword[200] ^ codeword[201] ^ codeword[203] ^ codeword[204] ^ codeword[206] ^ codeword[207] ^ codeword[210] ^ codeword[212] ^ codeword[213] ^ codeword[216] ^ codeword[219] ^ codeword[221] ^ codeword[222] ^ codeword[224] ^ codeword[225] ^ codeword[226] ^ codeword[228] ^ codeword[229] ^ codeword[231] ^ codeword[232] ^ codeword[235] ^ codeword[236] ^ codeword[238] ^ codeword[239] ^ codeword[241] ^ codeword[242] ^ codeword[245] ^ codeword[247] ^ codeword[248] ^ codeword[251] ^ codeword[254] ^ codeword[256] ^ codeword[258] ^ codeword[259] ^ codeword[261] ^ codeword[262] ^ codeword[265] ^ codeword[267] ^ codeword[268] ^ codeword[271] ^ codeword[274] ^ codeword[277] ^ codeword[278] ^ codeword[281] ^ codeword[284] ^ codeword[288] ^ codeword[291] ^ codeword[292] ^ codeword[294] ^ codeword[295] ^ codeword[296] ^ codeword[298] ^ codeword[299] ^ codeword[301] ^ codeword[302] ^ codeword[305] ^ codeword[306] ^ codeword[308] ^ codeword[309] ^ codeword[311] ^ codeword[312] ^ codeword[315] ^ codeword[317] ^ codeword[318] ^ codeword[321] ^ codeword[324] ^ codeword[326] ^ codeword[328] ^ codeword[329] ^ codeword[331] ^ codeword[332] ^ codeword[335] ^ codeword[337] ^ codeword[338] ^ codeword[341] ^ codeword[344] ^ codeword[347] ^ codeword[348] ^ codeword[351] ^ codeword[354] ^ codeword[358] ^ codeword[361] ^ codeword[363] ^ codeword[364] ^ codeword[366] ^ codeword[367] ^ codeword[370] ^ codeword[372] ^ codeword[373] ^ codeword[376] ^ codeword[379] ^ codeword[382] ^ codeword[383] ^ codeword[386] ^ codeword[389] ^ codeword[393] ^ codeword[397] ^ codeword[398] ^ codeword[401] ^ codeword[404] ^ codeword[408] ^ codeword[413] ^ codeword[417] ^ codeword[418] ^ codeword[420] ^ codeword[421] ^ codeword[422] ^ codeword[424] ^ codeword[425] ^ codeword[427] ^ codeword[428] ^ codeword[431] ^ codeword[432] ^ codeword[434] ^ codeword[435] ^ codeword[437] ^ codeword[438] ^ codeword[441] ^ codeword[443] ^ codeword[444] ^ codeword[447] ^ codeword[450] ^ codeword[452] ^ codeword[454] ^ codeword[455] ^ codeword[457] ^ codeword[458] ^ codeword[461] ^ codeword[463] ^ codeword[464] ^ codeword[467] ^ codeword[470] ^ codeword[473] ^ codeword[474] ^ codeword[477] ^ codeword[480] ^ codeword[484] ^ codeword[487] ^ codeword[489] ^ codeword[490] ^ codeword[492] ^ codeword[493] ^ codeword[496] ^ codeword[498] ^ codeword[499] ^ codeword[502] ^ codeword[505] ^ codeword[508] ^ codeword[509] ^ codeword[520];
    assign syndrome[9] = codeword[0] ^ codeword[1] ^ codeword[3] ^ codeword[4] ^ codeword[6] ^ codeword[8] ^ codeword[10] ^ codeword[12] ^ codeword[14] ^ codeword[17] ^ codeword[20] ^ codeword[22] ^ codeword[24] ^ codeword[27] ^ codeword[31] ^ codeword[35] ^ codeword[37] ^ codeword[39] ^ codeword[42] ^ codeword[46] ^ codeword[51] ^ codeword[56] ^ codeword[58] ^ codeword[60] ^ codeword[63] ^ codeword[67] ^ codeword[72] ^ codeword[78] ^ codeword[84] ^ codeword[86] ^ codeword[88] ^ codeword[91] ^ codeword[95] ^ codeword[100] ^ codeword[106] ^ codeword[113] ^ codeword[120] ^ codeword[122] ^ codeword[124] ^ codeword[127] ^ codeword[131] ^ codeword[136] ^ codeword[142] ^ codeword[149] ^ codeword[157] ^ codeword[165] ^ codeword[166] ^ codeword[167] ^ codeword[168] ^ codeword[170] ^ codeword[171] ^ codeword[172] ^ codeword[173] ^ codeword[175] ^ codeword[176] ^ codeword[177] ^ codeword[179] ^ codeword[180] ^ codeword[182] ^ codeword[184] ^ codeword[186] ^ codeword[187] ^ codeword[188] ^ codeword[190] ^ codeword[191] ^ codeword[192] ^ codeword[194] ^ codeword[195] ^ codeword[197] ^ codeword[199] ^ codeword[201] ^ codeword[202] ^ codeword[204] ^ codeword[205] ^ codeword[207] ^ codeword[209] ^ codeword[211] ^ codeword[213] ^ codeword[215] ^ codeword[218] ^ codeword[221] ^ codeword[222] ^ codeword[223] ^ codeword[225] ^ codeword[226] ^ codeword[227] ^ codeword[229] ^ codeword[230] ^ codeword[232] ^ codeword[234] ^ codeword[236] ^ codeword[237] ^ codeword[239] ^ codeword[240] ^ codeword[242] ^ codeword[244] ^ codeword[246] ^ codeword[248] ^ codeword[250] ^ codeword[253] ^ codeword[256] ^ codeword[257] ^ codeword[259] ^ codeword[260] ^ codeword[262] ^ codeword[264] ^ codeword[266] ^ codeword[268] ^ codeword[270] ^ codeword[273] ^ codeword[276] ^ codeword[278] ^ codeword[280] ^ codeword[283] ^ codeword[287] ^ codeword[291] ^ codeword[292] ^ codeword[293] ^ codeword[295] ^ codeword[296] ^ codeword[297] ^ codeword[299] ^ codeword[300] ^ codeword[302] ^ codeword[304] ^ codeword[306] ^ codeword[307] ^ codeword[309] ^ codeword[310] ^ codeword[312] ^ codeword[314] ^ codeword[316] ^ codeword[318] ^ codeword[320] ^ codeword[323] ^ codeword[326] ^ codeword[327] ^ codeword[329] ^ codeword[330] ^ codeword[332] ^ codeword[334] ^ codeword[336] ^ codeword[338] ^ codeword[340] ^ codeword[343] ^ codeword[346] ^ codeword[348] ^ codeword[350] ^ codeword[353] ^ codeword[357] ^ codeword[361] ^ codeword[362] ^ codeword[364] ^ codeword[365] ^ codeword[367] ^ codeword[369] ^ codeword[371] ^ codeword[373] ^ codeword[375] ^ codeword[378] ^ codeword[381] ^ codeword[383] ^ codeword[385] ^ codeword[388] ^ codeword[392] ^ codeword[396] ^ codeword[398] ^ codeword[400] ^ codeword[403] ^ codeword[407] ^ codeword[412] ^ codeword[417] ^ codeword[418] ^ codeword[419] ^ codeword[421] ^ codeword[422] ^ codeword[423] ^ codeword[425] ^ codeword[426] ^ codeword[428] ^ codeword[430] ^ codeword[432] ^ codeword[433] ^ codeword[435] ^ codeword[436] ^ codeword[438] ^ codeword[440] ^ codeword[442] ^ codeword[444] ^ codeword[446] ^ codeword[449] ^ codeword[452] ^ codeword[453] ^ codeword[455] ^ codeword[456] ^ codeword[458] ^ codeword[460] ^ codeword[462] ^ codeword[464] ^ codeword[466] ^ codeword[469] ^ codeword[472] ^ codeword[474] ^ codeword[476] ^ codeword[479] ^ codeword[483] ^ codeword[487] ^ codeword[488] ^ codeword[490] ^ codeword[491] ^ codeword[493] ^ codeword[495] ^ codeword[497] ^ codeword[499] ^ codeword[501] ^ codeword[504] ^ codeword[507] ^ codeword[509] ^ codeword[511] ^ codeword[521];
    assign syndrome[10] = codeword[0] ^ codeword[1] ^ codeword[2] ^ codeword[4] ^ codeword[5] ^ codeword[7] ^ codeword[10] ^ codeword[11] ^ codeword[13] ^ codeword[16] ^ codeword[20] ^ codeword[21] ^ codeword[23] ^ codeword[26] ^ codeword[30] ^ codeword[35] ^ codeword[36] ^ codeword[38] ^ codeword[41] ^ codeword[45] ^ codeword[50] ^ codeword[56] ^ codeword[57] ^ codeword[59] ^ codeword[62] ^ codeword[66] ^ codeword[71] ^ codeword[77] ^ codeword[84] ^ codeword[85] ^ codeword[87] ^ codeword[90] ^ codeword[94] ^ codeword[99] ^ codeword[105] ^ codeword[112] ^ codeword[120] ^ codeword[121] ^ codeword[123] ^ codeword[126] ^ codeword[130] ^ codeword[135] ^ codeword[141] ^ codeword[148] ^ codeword[156] ^ codeword[165] ^ codeword[166] ^ codeword[167] ^ codeword[168] ^ codeword[169] ^ codeword[171] ^ codeword[172] ^ codeword[173] ^ codeword[174] ^ codeword[176] ^ codeword[177] ^ codeword[178] ^ codeword[180] ^ codeword[181] ^ codeword[183] ^ codeword[186] ^ codeword[187] ^ codeword[188] ^ codeword[189] ^ codeword[191] ^ codeword[192] ^ codeword[193] ^ codeword[195] ^ codeword[196] ^ codeword[198] ^ codeword[201] ^ codeword[202] ^ codeword[203] ^ codeword[205] ^ codeword[206] ^ codeword[208] ^ codeword[211] ^ codeword[212] ^ codeword[214] ^ codeword[217] ^ codeword[221] ^ codeword[222] ^ codeword[223] ^ codeword[224] ^ codeword[226] ^ codeword[227] ^ codeword[228] ^ codeword[230] ^ codeword[231] ^ codeword[233] ^ codeword[236] ^ codeword[237] ^ codeword[238] ^ codeword[240] ^ codeword[241] ^ codeword[243] ^ codeword[246] ^ codeword[247] ^ codeword[249] ^ codeword[252] ^ codeword[256] ^ codeword[257] ^ codeword[258] ^ codeword[260] ^ codeword[261] ^ codeword[263] ^ codeword[266] ^ codeword[267] ^ codeword[269] ^ codeword[272] ^ codeword[276] ^ codeword[277] ^ codeword[279] ^ codeword[282] ^ codeword[286] ^ codeword[291] ^ codeword[292] ^ codeword[293] ^ codeword[294] ^ codeword[296] ^ codeword[297] ^ codeword[298] ^ codeword[300] ^ codeword[301] ^ codeword[303] ^ codeword[306] ^ codeword[307] ^ codeword[308] ^ codeword[310] ^ codeword[311] ^ codeword[313] ^ codeword[316] ^ codeword[317] ^ codeword[319] ^ codeword[322] ^ codeword[326] ^ codeword[327] ^ codeword[328] ^ codeword[330] ^ codeword[331] ^ codeword[333] ^ codeword[336] ^ codeword[337] ^ codeword[339] ^ codeword[342] ^ codeword[346] ^ codeword[347] ^ codeword[349] ^ codeword[352] ^ codeword[356] ^ codeword[361] ^ codeword[362] ^ codeword[363] ^ codeword[365] ^ codeword[366] ^ codeword[368] ^ codeword[371] ^ codeword[372] ^ codeword[374] ^ codeword[377] ^ codeword[381] ^ codeword[382] ^ codeword[384] ^ codeword[387] ^ codeword[391] ^ codeword[396] ^ codeword[397] ^ codeword[399] ^ codeword[402] ^ codeword[406] ^ codeword[411] ^ codeword[417] ^ codeword[418] ^ codeword[419] ^ codeword[420] ^ codeword[422] ^ codeword[423] ^ codeword[424] ^ codeword[426] ^ codeword[427] ^ codeword[429] ^ codeword[432] ^ codeword[433] ^ codeword[434] ^ codeword[436] ^ codeword[437] ^ codeword[439] ^ codeword[442] ^ codeword[443] ^ codeword[445] ^ codeword[448] ^ codeword[452] ^ codeword[453] ^ codeword[454] ^ codeword[456] ^ codeword[457] ^ codeword[459] ^ codeword[462] ^ codeword[463] ^ codeword[465] ^ codeword[468] ^ codeword[472] ^ codeword[473] ^ codeword[475] ^ codeword[478] ^ codeword[482] ^ codeword[487] ^ codeword[488] ^ codeword[489] ^ codeword[491] ^ codeword[492] ^ codeword[494] ^ codeword[497] ^ codeword[498] ^ codeword[500] ^ codeword[503] ^ codeword[507] ^ codeword[508] ^ codeword[510] ^ codeword[522];
  end else if (CodewordWidth == 1036 && MessageWidth == 1024) begin : gen_1036_1024
    `BR_ASSERT_STATIC(parity_width_matches_a, ParityWidth == 12)
    assign syndrome[0] = codeword[165] ^ codeword[166] ^ codeword[167] ^ codeword[168] ^ codeword[169] ^ codeword[170] ^ codeword[171] ^ codeword[172] ^ codeword[173] ^ codeword[174] ^ codeword[175] ^ codeword[176] ^ codeword[177] ^ codeword[178] ^ codeword[179] ^ codeword[180] ^ codeword[181] ^ codeword[182] ^ codeword[183] ^ codeword[184] ^ codeword[185] ^ codeword[186] ^ codeword[187] ^ codeword[188] ^ codeword[189] ^ codeword[190] ^ codeword[191] ^ codeword[192] ^ codeword[193] ^ codeword[194] ^ codeword[195] ^ codeword[196] ^ codeword[197] ^ codeword[198] ^ codeword[199] ^ codeword[200] ^ codeword[201] ^ codeword[202] ^ codeword[203] ^ codeword[204] ^ codeword[205] ^ codeword[206] ^ codeword[207] ^ codeword[208] ^ codeword[209] ^ codeword[210] ^ codeword[211] ^ codeword[212] ^ codeword[213] ^ codeword[214] ^ codeword[215] ^ codeword[216] ^ codeword[217] ^ codeword[218] ^ codeword[219] ^ codeword[682] ^ codeword[683] ^ codeword[684] ^ codeword[685] ^ codeword[686] ^ codeword[687] ^ codeword[688] ^ codeword[689] ^ codeword[690] ^ codeword[691] ^ codeword[692] ^ codeword[693] ^ codeword[694] ^ codeword[695] ^ codeword[696] ^ codeword[697] ^ codeword[698] ^ codeword[699] ^ codeword[700] ^ codeword[701] ^ codeword[702] ^ codeword[703] ^ codeword[704] ^ codeword[705] ^ codeword[706] ^ codeword[707] ^ codeword[708] ^ codeword[709] ^ codeword[710] ^ codeword[711] ^ codeword[712] ^ codeword[713] ^ codeword[714] ^ codeword[715] ^ codeword[716] ^ codeword[717] ^ codeword[718] ^ codeword[719] ^ codeword[720] ^ codeword[721] ^ codeword[722] ^ codeword[723] ^ codeword[724] ^ codeword[725] ^ codeword[726] ^ codeword[727] ^ codeword[728] ^ codeword[729] ^ codeword[730] ^ codeword[731] ^ codeword[732] ^ codeword[733] ^ codeword[734] ^ codeword[735] ^ codeword[736] ^ codeword[737] ^ codeword[738] ^ codeword[739] ^ codeword[740] ^ codeword[741] ^ codeword[742] ^ codeword[743] ^ codeword[744] ^ codeword[745] ^ codeword[746] ^ codeword[747] ^ codeword[748] ^ codeword[749] ^ codeword[750] ^ codeword[751] ^ codeword[752] ^ codeword[753] ^ codeword[754] ^ codeword[755] ^ codeword[756] ^ codeword[757] ^ codeword[758] ^ codeword[759] ^ codeword[760] ^ codeword[761] ^ codeword[762] ^ codeword[763] ^ codeword[764] ^ codeword[765] ^ codeword[766] ^ codeword[767] ^ codeword[768] ^ codeword[769] ^ codeword[770] ^ codeword[771] ^ codeword[772] ^ codeword[773] ^ codeword[774] ^ codeword[775] ^ codeword[776] ^ codeword[777] ^ codeword[778] ^ codeword[779] ^ codeword[780] ^ codeword[781] ^ codeword[782] ^ codeword[783] ^ codeword[784] ^ codeword[785] ^ codeword[786] ^ codeword[787] ^ codeword[788] ^ codeword[789] ^ codeword[790] ^ codeword[791] ^ codeword[792] ^ codeword[793] ^ codeword[794] ^ codeword[795] ^ codeword[796] ^ codeword[797] ^ codeword[798] ^ codeword[799] ^ codeword[800] ^ codeword[801] ^ codeword[802] ^ codeword[803] ^ codeword[804] ^ codeword[805] ^ codeword[806] ^ codeword[807] ^ codeword[808] ^ codeword[809] ^ codeword[810] ^ codeword[811] ^ codeword[812] ^ codeword[813] ^ codeword[814] ^ codeword[815] ^ codeword[816] ^ codeword[817] ^ codeword[818] ^ codeword[819] ^ codeword[820] ^ codeword[821] ^ codeword[822] ^ codeword[823] ^ codeword[824] ^ codeword[825] ^ codeword[826] ^ codeword[827] ^ codeword[828] ^ codeword[829] ^ codeword[830] ^ codeword[831] ^ codeword[832] ^ codeword[833] ^ codeword[834] ^ codeword[835] ^ codeword[836] ^ codeword[837] ^ codeword[838] ^ codeword[839] ^ codeword[840] ^ codeword[841] ^ codeword[842] ^ codeword[843] ^ codeword[844] ^ codeword[845] ^ codeword[846] ^ codeword[847] ^ codeword[848] ^ codeword[849] ^ codeword[850] ^ codeword[851] ^ codeword[852] ^ codeword[853] ^ codeword[854] ^ codeword[855] ^ codeword[856] ^ codeword[857] ^ codeword[858] ^ codeword[859] ^ codeword[860] ^ codeword[861] ^ codeword[862] ^ codeword[863] ^ codeword[864] ^ codeword[865] ^ codeword[866] ^ codeword[867] ^ codeword[868] ^ codeword[869] ^ codeword[870] ^ codeword[871] ^ codeword[872] ^ codeword[873] ^ codeword[874] ^ codeword[875] ^ codeword[876] ^ codeword[877] ^ codeword[878] ^ codeword[879] ^ codeword[880] ^ codeword[881] ^ codeword[882] ^ codeword[883] ^ codeword[884] ^ codeword[885] ^ codeword[886] ^ codeword[887] ^ codeword[888] ^ codeword[889] ^ codeword[890] ^ codeword[891] ^ codeword[892] ^ codeword[893] ^ codeword[894] ^ codeword[895] ^ codeword[896] ^ codeword[897] ^ codeword[898] ^ codeword[899] ^ codeword[900] ^ codeword[901] ^ codeword[902] ^ codeword[903] ^ codeword[904] ^ codeword[905] ^ codeword[906] ^ codeword[907] ^ codeword[908] ^ codeword[909] ^ codeword[910] ^ codeword[911] ^ codeword[912] ^ codeword[913] ^ codeword[914] ^ codeword[915] ^ codeword[916] ^ codeword[917] ^ codeword[918] ^ codeword[919] ^ codeword[920] ^ codeword[921] ^ codeword[922] ^ codeword[923] ^ codeword[924] ^ codeword[925] ^ codeword[926] ^ codeword[927] ^ codeword[928] ^ codeword[929] ^ codeword[930] ^ codeword[931] ^ codeword[932] ^ codeword[933] ^ codeword[934] ^ codeword[935] ^ codeword[936] ^ codeword[937] ^ codeword[938] ^ codeword[939] ^ codeword[940] ^ codeword[941] ^ codeword[942] ^ codeword[943] ^ codeword[944] ^ codeword[945] ^ codeword[946] ^ codeword[947] ^ codeword[948] ^ codeword[949] ^ codeword[950] ^ codeword[951] ^ codeword[952] ^ codeword[953] ^ codeword[954] ^ codeword[955] ^ codeword[956] ^ codeword[957] ^ codeword[958] ^ codeword[959] ^ codeword[960] ^ codeword[961] ^ codeword[962] ^ codeword[963] ^ codeword[964] ^ codeword[965] ^ codeword[966] ^ codeword[967] ^ codeword[968] ^ codeword[969] ^ codeword[970] ^ codeword[971] ^ codeword[972] ^ codeword[973] ^ codeword[974] ^ codeword[975] ^ codeword[976] ^ codeword[977] ^ codeword[978] ^ codeword[979] ^ codeword[980] ^ codeword[981] ^ codeword[982] ^ codeword[983] ^ codeword[984] ^ codeword[985] ^ codeword[986] ^ codeword[987] ^ codeword[988] ^ codeword[989] ^ codeword[990] ^ codeword[991] ^ codeword[992] ^ codeword[993] ^ codeword[994] ^ codeword[995] ^ codeword[996] ^ codeword[997] ^ codeword[998] ^ codeword[999] ^ codeword[1000] ^ codeword[1001] ^ codeword[1002] ^ codeword[1003] ^ codeword[1004] ^ codeword[1005] ^ codeword[1006] ^ codeword[1007] ^ codeword[1008] ^ codeword[1009] ^ codeword[1010] ^ codeword[1011] ^ codeword[1024];
    assign syndrome[1] = codeword[120] ^ codeword[121] ^ codeword[122] ^ codeword[123] ^ codeword[124] ^ codeword[125] ^ codeword[126] ^ codeword[127] ^ codeword[128] ^ codeword[129] ^ codeword[130] ^ codeword[131] ^ codeword[132] ^ codeword[133] ^ codeword[134] ^ codeword[135] ^ codeword[136] ^ codeword[137] ^ codeword[138] ^ codeword[139] ^ codeword[140] ^ codeword[141] ^ codeword[142] ^ codeword[143] ^ codeword[144] ^ codeword[145] ^ codeword[146] ^ codeword[147] ^ codeword[148] ^ codeword[149] ^ codeword[150] ^ codeword[151] ^ codeword[152] ^ codeword[153] ^ codeword[154] ^ codeword[155] ^ codeword[156] ^ codeword[157] ^ codeword[158] ^ codeword[159] ^ codeword[160] ^ codeword[161] ^ codeword[162] ^ codeword[163] ^ codeword[164] ^ codeword[210] ^ codeword[211] ^ codeword[212] ^ codeword[213] ^ codeword[214] ^ codeword[215] ^ codeword[216] ^ codeword[217] ^ codeword[218] ^ codeword[219] ^ codeword[472] ^ codeword[473] ^ codeword[474] ^ codeword[475] ^ codeword[476] ^ codeword[477] ^ codeword[478] ^ codeword[479] ^ codeword[480] ^ codeword[481] ^ codeword[482] ^ codeword[483] ^ codeword[484] ^ codeword[485] ^ codeword[486] ^ codeword[487] ^ codeword[488] ^ codeword[489] ^ codeword[490] ^ codeword[491] ^ codeword[492] ^ codeword[493] ^ codeword[494] ^ codeword[495] ^ codeword[496] ^ codeword[497] ^ codeword[498] ^ codeword[499] ^ codeword[500] ^ codeword[501] ^ codeword[502] ^ codeword[503] ^ codeword[504] ^ codeword[505] ^ codeword[506] ^ codeword[507] ^ codeword[508] ^ codeword[509] ^ codeword[510] ^ codeword[511] ^ codeword[512] ^ codeword[513] ^ codeword[514] ^ codeword[515] ^ codeword[516] ^ codeword[517] ^ codeword[518] ^ codeword[519] ^ codeword[520] ^ codeword[521] ^ codeword[522] ^ codeword[523] ^ codeword[524] ^ codeword[525] ^ codeword[526] ^ codeword[527] ^ codeword[528] ^ codeword[529] ^ codeword[530] ^ codeword[531] ^ codeword[532] ^ codeword[533] ^ codeword[534] ^ codeword[535] ^ codeword[536] ^ codeword[537] ^ codeword[538] ^ codeword[539] ^ codeword[540] ^ codeword[541] ^ codeword[542] ^ codeword[543] ^ codeword[544] ^ codeword[545] ^ codeword[546] ^ codeword[547] ^ codeword[548] ^ codeword[549] ^ codeword[550] ^ codeword[551] ^ codeword[552] ^ codeword[553] ^ codeword[554] ^ codeword[555] ^ codeword[556] ^ codeword[557] ^ codeword[558] ^ codeword[559] ^ codeword[560] ^ codeword[561] ^ codeword[562] ^ codeword[563] ^ codeword[564] ^ codeword[565] ^ codeword[566] ^ codeword[567] ^ codeword[568] ^ codeword[569] ^ codeword[570] ^ codeword[571] ^ codeword[572] ^ codeword[573] ^ codeword[574] ^ codeword[575] ^ codeword[576] ^ codeword[577] ^ codeword[578] ^ codeword[579] ^ codeword[580] ^ codeword[581] ^ codeword[582] ^ codeword[583] ^ codeword[584] ^ codeword[585] ^ codeword[586] ^ codeword[587] ^ codeword[588] ^ codeword[589] ^ codeword[590] ^ codeword[591] ^ codeword[592] ^ codeword[593] ^ codeword[594] ^ codeword[595] ^ codeword[596] ^ codeword[597] ^ codeword[598] ^ codeword[599] ^ codeword[600] ^ codeword[601] ^ codeword[602] ^ codeword[603] ^ codeword[604] ^ codeword[605] ^ codeword[606] ^ codeword[607] ^ codeword[608] ^ codeword[609] ^ codeword[610] ^ codeword[611] ^ codeword[612] ^ codeword[613] ^ codeword[614] ^ codeword[615] ^ codeword[616] ^ codeword[617] ^ codeword[618] ^ codeword[619] ^ codeword[620] ^ codeword[621] ^ codeword[622] ^ codeword[623] ^ codeword[624] ^ codeword[625] ^ codeword[626] ^ codeword[627] ^ codeword[628] ^ codeword[629] ^ codeword[630] ^ codeword[631] ^ codeword[632] ^ codeword[633] ^ codeword[634] ^ codeword[635] ^ codeword[636] ^ codeword[637] ^ codeword[638] ^ codeword[639] ^ codeword[640] ^ codeword[641] ^ codeword[642] ^ codeword[643] ^ codeword[644] ^ codeword[645] ^ codeword[646] ^ codeword[647] ^ codeword[648] ^ codeword[649] ^ codeword[650] ^ codeword[651] ^ codeword[652] ^ codeword[653] ^ codeword[654] ^ codeword[655] ^ codeword[656] ^ codeword[657] ^ codeword[658] ^ codeword[659] ^ codeword[660] ^ codeword[661] ^ codeword[662] ^ codeword[663] ^ codeword[664] ^ codeword[665] ^ codeword[666] ^ codeword[667] ^ codeword[668] ^ codeword[669] ^ codeword[670] ^ codeword[671] ^ codeword[672] ^ codeword[673] ^ codeword[674] ^ codeword[675] ^ codeword[676] ^ codeword[677] ^ codeword[678] ^ codeword[679] ^ codeword[680] ^ codeword[681] ^ codeword[892] ^ codeword[893] ^ codeword[894] ^ codeword[895] ^ codeword[896] ^ codeword[897] ^ codeword[898] ^ codeword[899] ^ codeword[900] ^ codeword[901] ^ codeword[902] ^ codeword[903] ^ codeword[904] ^ codeword[905] ^ codeword[906] ^ codeword[907] ^ codeword[908] ^ codeword[909] ^ codeword[910] ^ codeword[911] ^ codeword[912] ^ codeword[913] ^ codeword[914] ^ codeword[915] ^ codeword[916] ^ codeword[917] ^ codeword[918] ^ codeword[919] ^ codeword[920] ^ codeword[921] ^ codeword[922] ^ codeword[923] ^ codeword[924] ^ codeword[925] ^ codeword[926] ^ codeword[927] ^ codeword[928] ^ codeword[929] ^ codeword[930] ^ codeword[931] ^ codeword[932] ^ codeword[933] ^ codeword[934] ^ codeword[935] ^ codeword[936] ^ codeword[937] ^ codeword[938] ^ codeword[939] ^ codeword[940] ^ codeword[941] ^ codeword[942] ^ codeword[943] ^ codeword[944] ^ codeword[945] ^ codeword[946] ^ codeword[947] ^ codeword[948] ^ codeword[949] ^ codeword[950] ^ codeword[951] ^ codeword[952] ^ codeword[953] ^ codeword[954] ^ codeword[955] ^ codeword[956] ^ codeword[957] ^ codeword[958] ^ codeword[959] ^ codeword[960] ^ codeword[961] ^ codeword[962] ^ codeword[963] ^ codeword[964] ^ codeword[965] ^ codeword[966] ^ codeword[967] ^ codeword[968] ^ codeword[969] ^ codeword[970] ^ codeword[971] ^ codeword[972] ^ codeword[973] ^ codeword[974] ^ codeword[975] ^ codeword[976] ^ codeword[977] ^ codeword[978] ^ codeword[979] ^ codeword[980] ^ codeword[981] ^ codeword[982] ^ codeword[983] ^ codeword[984] ^ codeword[985] ^ codeword[986] ^ codeword[987] ^ codeword[988] ^ codeword[989] ^ codeword[990] ^ codeword[991] ^ codeword[992] ^ codeword[993] ^ codeword[994] ^ codeword[995] ^ codeword[996] ^ codeword[997] ^ codeword[998] ^ codeword[999] ^ codeword[1000] ^ codeword[1001] ^ codeword[1002] ^ codeword[1003] ^ codeword[1004] ^ codeword[1005] ^ codeword[1006] ^ codeword[1007] ^ codeword[1008] ^ codeword[1009] ^ codeword[1010] ^ codeword[1011] ^ codeword[1025];
    assign syndrome[2] = codeword[84] ^ codeword[85] ^ codeword[86] ^ codeword[87] ^ codeword[88] ^ codeword[89] ^ codeword[90] ^ codeword[91] ^ codeword[92] ^ codeword[93] ^ codeword[94] ^ codeword[95] ^ codeword[96] ^ codeword[97] ^ codeword[98] ^ codeword[99] ^ codeword[100] ^ codeword[101] ^ codeword[102] ^ codeword[103] ^ codeword[104] ^ codeword[105] ^ codeword[106] ^ codeword[107] ^ codeword[108] ^ codeword[109] ^ codeword[110] ^ codeword[111] ^ codeword[112] ^ codeword[113] ^ codeword[114] ^ codeword[115] ^ codeword[116] ^ codeword[117] ^ codeword[118] ^ codeword[119] ^ codeword[156] ^ codeword[157] ^ codeword[158] ^ codeword[159] ^ codeword[160] ^ codeword[161] ^ codeword[162] ^ codeword[163] ^ codeword[164] ^ codeword[201] ^ codeword[202] ^ codeword[203] ^ codeword[204] ^ codeword[205] ^ codeword[206] ^ codeword[207] ^ codeword[208] ^ codeword[209] ^ codeword[219] ^ codeword[346] ^ codeword[347] ^ codeword[348] ^ codeword[349] ^ codeword[350] ^ codeword[351] ^ codeword[352] ^ codeword[353] ^ codeword[354] ^ codeword[355] ^ codeword[356] ^ codeword[357] ^ codeword[358] ^ codeword[359] ^ codeword[360] ^ codeword[361] ^ codeword[362] ^ codeword[363] ^ codeword[364] ^ codeword[365] ^ codeword[366] ^ codeword[367] ^ codeword[368] ^ codeword[369] ^ codeword[370] ^ codeword[371] ^ codeword[372] ^ codeword[373] ^ codeword[374] ^ codeword[375] ^ codeword[376] ^ codeword[377] ^ codeword[378] ^ codeword[379] ^ codeword[380] ^ codeword[381] ^ codeword[382] ^ codeword[383] ^ codeword[384] ^ codeword[385] ^ codeword[386] ^ codeword[387] ^ codeword[388] ^ codeword[389] ^ codeword[390] ^ codeword[391] ^ codeword[392] ^ codeword[393] ^ codeword[394] ^ codeword[395] ^ codeword[396] ^ codeword[397] ^ codeword[398] ^ codeword[399] ^ codeword[400] ^ codeword[401] ^ codeword[402] ^ codeword[403] ^ codeword[404] ^ codeword[405] ^ codeword[406] ^ codeword[407] ^ codeword[408] ^ codeword[409] ^ codeword[410] ^ codeword[411] ^ codeword[412] ^ codeword[413] ^ codeword[414] ^ codeword[415] ^ codeword[416] ^ codeword[417] ^ codeword[418] ^ codeword[419] ^ codeword[420] ^ codeword[421] ^ codeword[422] ^ codeword[423] ^ codeword[424] ^ codeword[425] ^ codeword[426] ^ codeword[427] ^ codeword[428] ^ codeword[429] ^ codeword[430] ^ codeword[431] ^ codeword[432] ^ codeword[433] ^ codeword[434] ^ codeword[435] ^ codeword[436] ^ codeword[437] ^ codeword[438] ^ codeword[439] ^ codeword[440] ^ codeword[441] ^ codeword[442] ^ codeword[443] ^ codeword[444] ^ codeword[445] ^ codeword[446] ^ codeword[447] ^ codeword[448] ^ codeword[449] ^ codeword[450] ^ codeword[451] ^ codeword[452] ^ codeword[453] ^ codeword[454] ^ codeword[455] ^ codeword[456] ^ codeword[457] ^ codeword[458] ^ codeword[459] ^ codeword[460] ^ codeword[461] ^ codeword[462] ^ codeword[463] ^ codeword[464] ^ codeword[465] ^ codeword[466] ^ codeword[467] ^ codeword[468] ^ codeword[469] ^ codeword[470] ^ codeword[471] ^ codeword[598] ^ codeword[599] ^ codeword[600] ^ codeword[601] ^ codeword[602] ^ codeword[603] ^ codeword[604] ^ codeword[605] ^ codeword[606] ^ codeword[607] ^ codeword[608] ^ codeword[609] ^ codeword[610] ^ codeword[611] ^ codeword[612] ^ codeword[613] ^ codeword[614] ^ codeword[615] ^ codeword[616] ^ codeword[617] ^ codeword[618] ^ codeword[619] ^ codeword[620] ^ codeword[621] ^ codeword[622] ^ codeword[623] ^ codeword[624] ^ codeword[625] ^ codeword[626] ^ codeword[627] ^ codeword[628] ^ codeword[629] ^ codeword[630] ^ codeword[631] ^ codeword[632] ^ codeword[633] ^ codeword[634] ^ codeword[635] ^ codeword[636] ^ codeword[637] ^ codeword[638] ^ codeword[639] ^ codeword[640] ^ codeword[641] ^ codeword[642] ^ codeword[643] ^ codeword[644] ^ codeword[645] ^ codeword[646] ^ codeword[647] ^ codeword[648] ^ codeword[649] ^ codeword[650] ^ codeword[651] ^ codeword[652] ^ codeword[653] ^ codeword[654] ^ codeword[655] ^ codeword[656] ^ codeword[657] ^ codeword[658] ^ codeword[659] ^ codeword[660] ^ codeword[661] ^ codeword[662] ^ codeword[663] ^ codeword[664] ^ codeword[665] ^ codeword[666] ^ codeword[667] ^ codeword[668] ^ codeword[669] ^ codeword[670] ^ codeword[671] ^ codeword[672] ^ codeword[673] ^ codeword[674] ^ codeword[675] ^ codeword[676] ^ codeword[677] ^ codeword[678] ^ codeword[679] ^ codeword[680] ^ codeword[681] ^ codeword[808] ^ codeword[809] ^ codeword[810] ^ codeword[811] ^ codeword[812] ^ codeword[813] ^ codeword[814] ^ codeword[815] ^ codeword[816] ^ codeword[817] ^ codeword[818] ^ codeword[819] ^ codeword[820] ^ codeword[821] ^ codeword[822] ^ codeword[823] ^ codeword[824] ^ codeword[825] ^ codeword[826] ^ codeword[827] ^ codeword[828] ^ codeword[829] ^ codeword[830] ^ codeword[831] ^ codeword[832] ^ codeword[833] ^ codeword[834] ^ codeword[835] ^ codeword[836] ^ codeword[837] ^ codeword[838] ^ codeword[839] ^ codeword[840] ^ codeword[841] ^ codeword[842] ^ codeword[843] ^ codeword[844] ^ codeword[845] ^ codeword[846] ^ codeword[847] ^ codeword[848] ^ codeword[849] ^ codeword[850] ^ codeword[851] ^ codeword[852] ^ codeword[853] ^ codeword[854] ^ codeword[855] ^ codeword[856] ^ codeword[857] ^ codeword[858] ^ codeword[859] ^ codeword[860] ^ codeword[861] ^ codeword[862] ^ codeword[863] ^ codeword[864] ^ codeword[865] ^ codeword[866] ^ codeword[867] ^ codeword[868] ^ codeword[869] ^ codeword[870] ^ codeword[871] ^ codeword[872] ^ codeword[873] ^ codeword[874] ^ codeword[875] ^ codeword[876] ^ codeword[877] ^ codeword[878] ^ codeword[879] ^ codeword[880] ^ codeword[881] ^ codeword[882] ^ codeword[883] ^ codeword[884] ^ codeword[885] ^ codeword[886] ^ codeword[887] ^ codeword[888] ^ codeword[889] ^ codeword[890] ^ codeword[891] ^ codeword[976] ^ codeword[977] ^ codeword[978] ^ codeword[979] ^ codeword[980] ^ codeword[981] ^ codeword[982] ^ codeword[983] ^ codeword[984] ^ codeword[985] ^ codeword[986] ^ codeword[987] ^ codeword[988] ^ codeword[989] ^ codeword[990] ^ codeword[991] ^ codeword[992] ^ codeword[993] ^ codeword[994] ^ codeword[995] ^ codeword[996] ^ codeword[997] ^ codeword[998] ^ codeword[999] ^ codeword[1000] ^ codeword[1001] ^ codeword[1002] ^ codeword[1003] ^ codeword[1004] ^ codeword[1005] ^ codeword[1006] ^ codeword[1007] ^ codeword[1008] ^ codeword[1009] ^ codeword[1010] ^ codeword[1011] ^ codeword[1026];
    assign syndrome[3] = codeword[56] ^ codeword[57] ^ codeword[58] ^ codeword[59] ^ codeword[60] ^ codeword[61] ^ codeword[62] ^ codeword[63] ^ codeword[64] ^ codeword[65] ^ codeword[66] ^ codeword[67] ^ codeword[68] ^ codeword[69] ^ codeword[70] ^ codeword[71] ^ codeword[72] ^ codeword[73] ^ codeword[74] ^ codeword[75] ^ codeword[76] ^ codeword[77] ^ codeword[78] ^ codeword[79] ^ codeword[80] ^ codeword[81] ^ codeword[82] ^ codeword[83] ^ codeword[112] ^ codeword[113] ^ codeword[114] ^ codeword[115] ^ codeword[116] ^ codeword[117] ^ codeword[118] ^ codeword[119] ^ codeword[148] ^ codeword[149] ^ codeword[150] ^ codeword[151] ^ codeword[152] ^ codeword[153] ^ codeword[154] ^ codeword[155] ^ codeword[164] ^ codeword[193] ^ codeword[194] ^ codeword[195] ^ codeword[196] ^ codeword[197] ^ codeword[198] ^ codeword[199] ^ codeword[200] ^ codeword[209] ^ codeword[218] ^ codeword[276] ^ codeword[277] ^ codeword[278] ^ codeword[279] ^ codeword[280] ^ codeword[281] ^ codeword[282] ^ codeword[283] ^ codeword[284] ^ codeword[285] ^ codeword[286] ^ codeword[287] ^ codeword[288] ^ codeword[289] ^ codeword[290] ^ codeword[291] ^ codeword[292] ^ codeword[293] ^ codeword[294] ^ codeword[295] ^ codeword[296] ^ codeword[297] ^ codeword[298] ^ codeword[299] ^ codeword[300] ^ codeword[301] ^ codeword[302] ^ codeword[303] ^ codeword[304] ^ codeword[305] ^ codeword[306] ^ codeword[307] ^ codeword[308] ^ codeword[309] ^ codeword[310] ^ codeword[311] ^ codeword[312] ^ codeword[313] ^ codeword[314] ^ codeword[315] ^ codeword[316] ^ codeword[317] ^ codeword[318] ^ codeword[319] ^ codeword[320] ^ codeword[321] ^ codeword[322] ^ codeword[323] ^ codeword[324] ^ codeword[325] ^ codeword[326] ^ codeword[327] ^ codeword[328] ^ codeword[329] ^ codeword[330] ^ codeword[331] ^ codeword[332] ^ codeword[333] ^ codeword[334] ^ codeword[335] ^ codeword[336] ^ codeword[337] ^ codeword[338] ^ codeword[339] ^ codeword[340] ^ codeword[341] ^ codeword[342] ^ codeword[343] ^ codeword[344] ^ codeword[345] ^ codeword[416] ^ codeword[417] ^ codeword[418] ^ codeword[419] ^ codeword[420] ^ codeword[421] ^ codeword[422] ^ codeword[423] ^ codeword[424] ^ codeword[425] ^ codeword[426] ^ codeword[427] ^ codeword[428] ^ codeword[429] ^ codeword[430] ^ codeword[431] ^ codeword[432] ^ codeword[433] ^ codeword[434] ^ codeword[435] ^ codeword[436] ^ codeword[437] ^ codeword[438] ^ codeword[439] ^ codeword[440] ^ codeword[441] ^ codeword[442] ^ codeword[443] ^ codeword[444] ^ codeword[445] ^ codeword[446] ^ codeword[447] ^ codeword[448] ^ codeword[449] ^ codeword[450] ^ codeword[451] ^ codeword[452] ^ codeword[453] ^ codeword[454] ^ codeword[455] ^ codeword[456] ^ codeword[457] ^ codeword[458] ^ codeword[459] ^ codeword[460] ^ codeword[461] ^ codeword[462] ^ codeword[463] ^ codeword[464] ^ codeword[465] ^ codeword[466] ^ codeword[467] ^ codeword[468] ^ codeword[469] ^ codeword[470] ^ codeword[471] ^ codeword[542] ^ codeword[543] ^ codeword[544] ^ codeword[545] ^ codeword[546] ^ codeword[547] ^ codeword[548] ^ codeword[549] ^ codeword[550] ^ codeword[551] ^ codeword[552] ^ codeword[553] ^ codeword[554] ^ codeword[555] ^ codeword[556] ^ codeword[557] ^ codeword[558] ^ codeword[559] ^ codeword[560] ^ codeword[561] ^ codeword[562] ^ codeword[563] ^ codeword[564] ^ codeword[565] ^ codeword[566] ^ codeword[567] ^ codeword[568] ^ codeword[569] ^ codeword[570] ^ codeword[571] ^ codeword[572] ^ codeword[573] ^ codeword[574] ^ codeword[575] ^ codeword[576] ^ codeword[577] ^ codeword[578] ^ codeword[579] ^ codeword[580] ^ codeword[581] ^ codeword[582] ^ codeword[583] ^ codeword[584] ^ codeword[585] ^ codeword[586] ^ codeword[587] ^ codeword[588] ^ codeword[589] ^ codeword[590] ^ codeword[591] ^ codeword[592] ^ codeword[593] ^ codeword[594] ^ codeword[595] ^ codeword[596] ^ codeword[597] ^ codeword[654] ^ codeword[655] ^ codeword[656] ^ codeword[657] ^ codeword[658] ^ codeword[659] ^ codeword[660] ^ codeword[661] ^ codeword[662] ^ codeword[663] ^ codeword[664] ^ codeword[665] ^ codeword[666] ^ codeword[667] ^ codeword[668] ^ codeword[669] ^ codeword[670] ^ codeword[671] ^ codeword[672] ^ codeword[673] ^ codeword[674] ^ codeword[675] ^ codeword[676] ^ codeword[677] ^ codeword[678] ^ codeword[679] ^ codeword[680] ^ codeword[681] ^ codeword[752] ^ codeword[753] ^ codeword[754] ^ codeword[755] ^ codeword[756] ^ codeword[757] ^ codeword[758] ^ codeword[759] ^ codeword[760] ^ codeword[761] ^ codeword[762] ^ codeword[763] ^ codeword[764] ^ codeword[765] ^ codeword[766] ^ codeword[767] ^ codeword[768] ^ codeword[769] ^ codeword[770] ^ codeword[771] ^ codeword[772] ^ codeword[773] ^ codeword[774] ^ codeword[775] ^ codeword[776] ^ codeword[777] ^ codeword[778] ^ codeword[779] ^ codeword[780] ^ codeword[781] ^ codeword[782] ^ codeword[783] ^ codeword[784] ^ codeword[785] ^ codeword[786] ^ codeword[787] ^ codeword[788] ^ codeword[789] ^ codeword[790] ^ codeword[791] ^ codeword[792] ^ codeword[793] ^ codeword[794] ^ codeword[795] ^ codeword[796] ^ codeword[797] ^ codeword[798] ^ codeword[799] ^ codeword[800] ^ codeword[801] ^ codeword[802] ^ codeword[803] ^ codeword[804] ^ codeword[805] ^ codeword[806] ^ codeword[807] ^ codeword[864] ^ codeword[865] ^ codeword[866] ^ codeword[867] ^ codeword[868] ^ codeword[869] ^ codeword[870] ^ codeword[871] ^ codeword[872] ^ codeword[873] ^ codeword[874] ^ codeword[875] ^ codeword[876] ^ codeword[877] ^ codeword[878] ^ codeword[879] ^ codeword[880] ^ codeword[881] ^ codeword[882] ^ codeword[883] ^ codeword[884] ^ codeword[885] ^ codeword[886] ^ codeword[887] ^ codeword[888] ^ codeword[889] ^ codeword[890] ^ codeword[891] ^ codeword[948] ^ codeword[949] ^ codeword[950] ^ codeword[951] ^ codeword[952] ^ codeword[953] ^ codeword[954] ^ codeword[955] ^ codeword[956] ^ codeword[957] ^ codeword[958] ^ codeword[959] ^ codeword[960] ^ codeword[961] ^ codeword[962] ^ codeword[963] ^ codeword[964] ^ codeword[965] ^ codeword[966] ^ codeword[967] ^ codeword[968] ^ codeword[969] ^ codeword[970] ^ codeword[971] ^ codeword[972] ^ codeword[973] ^ codeword[974] ^ codeword[975] ^ codeword[1004] ^ codeword[1005] ^ codeword[1006] ^ codeword[1007] ^ codeword[1008] ^ codeword[1009] ^ codeword[1010] ^ codeword[1011] ^ codeword[1020] ^ codeword[1021] ^ codeword[1022] ^ codeword[1023] ^ codeword[1027];
    assign syndrome[4] = codeword[35] ^ codeword[36] ^ codeword[37] ^ codeword[38] ^ codeword[39] ^ codeword[40] ^ codeword[41] ^ codeword[42] ^ codeword[43] ^ codeword[44] ^ codeword[45] ^ codeword[46] ^ codeword[47] ^ codeword[48] ^ codeword[49] ^ codeword[50] ^ codeword[51] ^ codeword[52] ^ codeword[53] ^ codeword[54] ^ codeword[55] ^ codeword[77] ^ codeword[78] ^ codeword[79] ^ codeword[80] ^ codeword[81] ^ codeword[82] ^ codeword[83] ^ codeword[105] ^ codeword[106] ^ codeword[107] ^ codeword[108] ^ codeword[109] ^ codeword[110] ^ codeword[111] ^ codeword[119] ^ codeword[141] ^ codeword[142] ^ codeword[143] ^ codeword[144] ^ codeword[145] ^ codeword[146] ^ codeword[147] ^ codeword[155] ^ codeword[163] ^ codeword[186] ^ codeword[187] ^ codeword[188] ^ codeword[189] ^ codeword[190] ^ codeword[191] ^ codeword[192] ^ codeword[200] ^ codeword[208] ^ codeword[217] ^ codeword[241] ^ codeword[242] ^ codeword[243] ^ codeword[244] ^ codeword[245] ^ codeword[246] ^ codeword[247] ^ codeword[248] ^ codeword[249] ^ codeword[250] ^ codeword[251] ^ codeword[252] ^ codeword[253] ^ codeword[254] ^ codeword[255] ^ codeword[256] ^ codeword[257] ^ codeword[258] ^ codeword[259] ^ codeword[260] ^ codeword[261] ^ codeword[262] ^ codeword[263] ^ codeword[264] ^ codeword[265] ^ codeword[266] ^ codeword[267] ^ codeword[268] ^ codeword[269] ^ codeword[270] ^ codeword[271] ^ codeword[272] ^ codeword[273] ^ codeword[274] ^ codeword[275] ^ codeword[311] ^ codeword[312] ^ codeword[313] ^ codeword[314] ^ codeword[315] ^ codeword[316] ^ codeword[317] ^ codeword[318] ^ codeword[319] ^ codeword[320] ^ codeword[321] ^ codeword[322] ^ codeword[323] ^ codeword[324] ^ codeword[325] ^ codeword[326] ^ codeword[327] ^ codeword[328] ^ codeword[329] ^ codeword[330] ^ codeword[331] ^ codeword[332] ^ codeword[333] ^ codeword[334] ^ codeword[335] ^ codeword[336] ^ codeword[337] ^ codeword[338] ^ codeword[339] ^ codeword[340] ^ codeword[341] ^ codeword[342] ^ codeword[343] ^ codeword[344] ^ codeword[345] ^ codeword[381] ^ codeword[382] ^ codeword[383] ^ codeword[384] ^ codeword[385] ^ codeword[386] ^ codeword[387] ^ codeword[388] ^ codeword[389] ^ codeword[390] ^ codeword[391] ^ codeword[392] ^ codeword[393] ^ codeword[394] ^ codeword[395] ^ codeword[396] ^ codeword[397] ^ codeword[398] ^ codeword[399] ^ codeword[400] ^ codeword[401] ^ codeword[402] ^ codeword[403] ^ codeword[404] ^ codeword[405] ^ codeword[406] ^ codeword[407] ^ codeword[408] ^ codeword[409] ^ codeword[410] ^ codeword[411] ^ codeword[412] ^ codeword[413] ^ codeword[414] ^ codeword[415] ^ codeword[451] ^ codeword[452] ^ codeword[453] ^ codeword[454] ^ codeword[455] ^ codeword[456] ^ codeword[457] ^ codeword[458] ^ codeword[459] ^ codeword[460] ^ codeword[461] ^ codeword[462] ^ codeword[463] ^ codeword[464] ^ codeword[465] ^ codeword[466] ^ codeword[467] ^ codeword[468] ^ codeword[469] ^ codeword[470] ^ codeword[471] ^ codeword[507] ^ codeword[508] ^ codeword[509] ^ codeword[510] ^ codeword[511] ^ codeword[512] ^ codeword[513] ^ codeword[514] ^ codeword[515] ^ codeword[516] ^ codeword[517] ^ codeword[518] ^ codeword[519] ^ codeword[520] ^ codeword[521] ^ codeword[522] ^ codeword[523] ^ codeword[524] ^ codeword[525] ^ codeword[526] ^ codeword[527] ^ codeword[528] ^ codeword[529] ^ codeword[530] ^ codeword[531] ^ codeword[532] ^ codeword[533] ^ codeword[534] ^ codeword[535] ^ codeword[536] ^ codeword[537] ^ codeword[538] ^ codeword[539] ^ codeword[540] ^ codeword[541] ^ codeword[577] ^ codeword[578] ^ codeword[579] ^ codeword[580] ^ codeword[581] ^ codeword[582] ^ codeword[583] ^ codeword[584] ^ codeword[585] ^ codeword[586] ^ codeword[587] ^ codeword[588] ^ codeword[589] ^ codeword[590] ^ codeword[591] ^ codeword[592] ^ codeword[593] ^ codeword[594] ^ codeword[595] ^ codeword[596] ^ codeword[597] ^ codeword[633] ^ codeword[634] ^ codeword[635] ^ codeword[636] ^ codeword[637] ^ codeword[638] ^ codeword[639] ^ codeword[640] ^ codeword[641] ^ codeword[642] ^ codeword[643] ^ codeword[644] ^ codeword[645] ^ codeword[646] ^ codeword[647] ^ codeword[648] ^ codeword[649] ^ codeword[650] ^ codeword[651] ^ codeword[652] ^ codeword[653] ^ codeword[675] ^ codeword[676] ^ codeword[677] ^ codeword[678] ^ codeword[679] ^ codeword[680] ^ codeword[681] ^ codeword[717] ^ codeword[718] ^ codeword[719] ^ codeword[720] ^ codeword[721] ^ codeword[722] ^ codeword[723] ^ codeword[724] ^ codeword[725] ^ codeword[726] ^ codeword[727] ^ codeword[728] ^ codeword[729] ^ codeword[730] ^ codeword[731] ^ codeword[732] ^ codeword[733] ^ codeword[734] ^ codeword[735] ^ codeword[736] ^ codeword[737] ^ codeword[738] ^ codeword[739] ^ codeword[740] ^ codeword[741] ^ codeword[742] ^ codeword[743] ^ codeword[744] ^ codeword[745] ^ codeword[746] ^ codeword[747] ^ codeword[748] ^ codeword[749] ^ codeword[750] ^ codeword[751] ^ codeword[787] ^ codeword[788] ^ codeword[789] ^ codeword[790] ^ codeword[791] ^ codeword[792] ^ codeword[793] ^ codeword[794] ^ codeword[795] ^ codeword[796] ^ codeword[797] ^ codeword[798] ^ codeword[799] ^ codeword[800] ^ codeword[801] ^ codeword[802] ^ codeword[803] ^ codeword[804] ^ codeword[805] ^ codeword[806] ^ codeword[807] ^ codeword[843] ^ codeword[844] ^ codeword[845] ^ codeword[846] ^ codeword[847] ^ codeword[848] ^ codeword[849] ^ codeword[850] ^ codeword[851] ^ codeword[852] ^ codeword[853] ^ codeword[854] ^ codeword[855] ^ codeword[856] ^ codeword[857] ^ codeword[858] ^ codeword[859] ^ codeword[860] ^ codeword[861] ^ codeword[862] ^ codeword[863] ^ codeword[885] ^ codeword[886] ^ codeword[887] ^ codeword[888] ^ codeword[889] ^ codeword[890] ^ codeword[891] ^ codeword[927] ^ codeword[928] ^ codeword[929] ^ codeword[930] ^ codeword[931] ^ codeword[932] ^ codeword[933] ^ codeword[934] ^ codeword[935] ^ codeword[936] ^ codeword[937] ^ codeword[938] ^ codeword[939] ^ codeword[940] ^ codeword[941] ^ codeword[942] ^ codeword[943] ^ codeword[944] ^ codeword[945] ^ codeword[946] ^ codeword[947] ^ codeword[969] ^ codeword[970] ^ codeword[971] ^ codeword[972] ^ codeword[973] ^ codeword[974] ^ codeword[975] ^ codeword[997] ^ codeword[998] ^ codeword[999] ^ codeword[1000] ^ codeword[1001] ^ codeword[1002] ^ codeword[1003] ^ codeword[1011] ^ codeword[1013] ^ codeword[1014] ^ codeword[1015] ^ codeword[1016] ^ codeword[1017] ^ codeword[1018] ^ codeword[1019] ^ codeword[1028];
    assign syndrome[5] = codeword[20] ^ codeword[21] ^ codeword[22] ^ codeword[23] ^ codeword[24] ^ codeword[25] ^ codeword[26] ^ codeword[27] ^ codeword[28] ^ codeword[29] ^ codeword[30] ^ codeword[31] ^ codeword[32] ^ codeword[33] ^ codeword[34] ^ codeword[50] ^ codeword[51] ^ codeword[52] ^ codeword[53] ^ codeword[54] ^ codeword[55] ^ codeword[71] ^ codeword[72] ^ codeword[73] ^ codeword[74] ^ codeword[75] ^ codeword[76] ^ codeword[83] ^ codeword[99] ^ codeword[100] ^ codeword[101] ^ codeword[102] ^ codeword[103] ^ codeword[104] ^ codeword[111] ^ codeword[118] ^ codeword[135] ^ codeword[136] ^ codeword[137] ^ codeword[138] ^ codeword[139] ^ codeword[140] ^ codeword[147] ^ codeword[154] ^ codeword[162] ^ codeword[180] ^ codeword[181] ^ codeword[182] ^ codeword[183] ^ codeword[184] ^ codeword[185] ^ codeword[192] ^ codeword[199] ^ codeword[207] ^ codeword[216] ^ codeword[226] ^ codeword[227] ^ codeword[228] ^ codeword[229] ^ codeword[230] ^ codeword[231] ^ codeword[232] ^ codeword[233] ^ codeword[234] ^ codeword[235] ^ codeword[236] ^ codeword[237] ^ codeword[238] ^ codeword[239] ^ codeword[240] ^ codeword[256] ^ codeword[257] ^ codeword[258] ^ codeword[259] ^ codeword[260] ^ codeword[261] ^ codeword[262] ^ codeword[263] ^ codeword[264] ^ codeword[265] ^ codeword[266] ^ codeword[267] ^ codeword[268] ^ codeword[269] ^ codeword[270] ^ codeword[271] ^ codeword[272] ^ codeword[273] ^ codeword[274] ^ codeword[275] ^ codeword[291] ^ codeword[292] ^ codeword[293] ^ codeword[294] ^ codeword[295] ^ codeword[296] ^ codeword[297] ^ codeword[298] ^ codeword[299] ^ codeword[300] ^ codeword[301] ^ codeword[302] ^ codeword[303] ^ codeword[304] ^ codeword[305] ^ codeword[306] ^ codeword[307] ^ codeword[308] ^ codeword[309] ^ codeword[310] ^ codeword[331] ^ codeword[332] ^ codeword[333] ^ codeword[334] ^ codeword[335] ^ codeword[336] ^ codeword[337] ^ codeword[338] ^ codeword[339] ^ codeword[340] ^ codeword[341] ^ codeword[342] ^ codeword[343] ^ codeword[344] ^ codeword[345] ^ codeword[361] ^ codeword[362] ^ codeword[363] ^ codeword[364] ^ codeword[365] ^ codeword[366] ^ codeword[367] ^ codeword[368] ^ codeword[369] ^ codeword[370] ^ codeword[371] ^ codeword[372] ^ codeword[373] ^ codeword[374] ^ codeword[375] ^ codeword[376] ^ codeword[377] ^ codeword[378] ^ codeword[379] ^ codeword[380] ^ codeword[401] ^ codeword[402] ^ codeword[403] ^ codeword[404] ^ codeword[405] ^ codeword[406] ^ codeword[407] ^ codeword[408] ^ codeword[409] ^ codeword[410] ^ codeword[411] ^ codeword[412] ^ codeword[413] ^ codeword[414] ^ codeword[415] ^ codeword[436] ^ codeword[437] ^ codeword[438] ^ codeword[439] ^ codeword[440] ^ codeword[441] ^ codeword[442] ^ codeword[443] ^ codeword[444] ^ codeword[445] ^ codeword[446] ^ codeword[447] ^ codeword[448] ^ codeword[449] ^ codeword[450] ^ codeword[466] ^ codeword[467] ^ codeword[468] ^ codeword[469] ^ codeword[470] ^ codeword[471] ^ codeword[487] ^ codeword[488] ^ codeword[489] ^ codeword[490] ^ codeword[491] ^ codeword[492] ^ codeword[493] ^ codeword[494] ^ codeword[495] ^ codeword[496] ^ codeword[497] ^ codeword[498] ^ codeword[499] ^ codeword[500] ^ codeword[501] ^ codeword[502] ^ codeword[503] ^ codeword[504] ^ codeword[505] ^ codeword[506] ^ codeword[527] ^ codeword[528] ^ codeword[529] ^ codeword[530] ^ codeword[531] ^ codeword[532] ^ codeword[533] ^ codeword[534] ^ codeword[535] ^ codeword[536] ^ codeword[537] ^ codeword[538] ^ codeword[539] ^ codeword[540] ^ codeword[541] ^ codeword[562] ^ codeword[563] ^ codeword[564] ^ codeword[565] ^ codeword[566] ^ codeword[567] ^ codeword[568] ^ codeword[569] ^ codeword[570] ^ codeword[571] ^ codeword[572] ^ codeword[573] ^ codeword[574] ^ codeword[575] ^ codeword[576] ^ codeword[592] ^ codeword[593] ^ codeword[594] ^ codeword[595] ^ codeword[596] ^ codeword[597] ^ codeword[618] ^ codeword[619] ^ codeword[620] ^ codeword[621] ^ codeword[622] ^ codeword[623] ^ codeword[624] ^ codeword[625] ^ codeword[626] ^ codeword[627] ^ codeword[628] ^ codeword[629] ^ codeword[630] ^ codeword[631] ^ codeword[632] ^ codeword[648] ^ codeword[649] ^ codeword[650] ^ codeword[651] ^ codeword[652] ^ codeword[653] ^ codeword[669] ^ codeword[670] ^ codeword[671] ^ codeword[672] ^ codeword[673] ^ codeword[674] ^ codeword[681] ^ codeword[697] ^ codeword[698] ^ codeword[699] ^ codeword[700] ^ codeword[701] ^ codeword[702] ^ codeword[703] ^ codeword[704] ^ codeword[705] ^ codeword[706] ^ codeword[707] ^ codeword[708] ^ codeword[709] ^ codeword[710] ^ codeword[711] ^ codeword[712] ^ codeword[713] ^ codeword[714] ^ codeword[715] ^ codeword[716] ^ codeword[737] ^ codeword[738] ^ codeword[739] ^ codeword[740] ^ codeword[741] ^ codeword[742] ^ codeword[743] ^ codeword[744] ^ codeword[745] ^ codeword[746] ^ codeword[747] ^ codeword[748] ^ codeword[749] ^ codeword[750] ^ codeword[751] ^ codeword[772] ^ codeword[773] ^ codeword[774] ^ codeword[775] ^ codeword[776] ^ codeword[777] ^ codeword[778] ^ codeword[779] ^ codeword[780] ^ codeword[781] ^ codeword[782] ^ codeword[783] ^ codeword[784] ^ codeword[785] ^ codeword[786] ^ codeword[802] ^ codeword[803] ^ codeword[804] ^ codeword[805] ^ codeword[806] ^ codeword[807] ^ codeword[828] ^ codeword[829] ^ codeword[830] ^ codeword[831] ^ codeword[832] ^ codeword[833] ^ codeword[834] ^ codeword[835] ^ codeword[836] ^ codeword[837] ^ codeword[838] ^ codeword[839] ^ codeword[840] ^ codeword[841] ^ codeword[842] ^ codeword[858] ^ codeword[859] ^ codeword[860] ^ codeword[861] ^ codeword[862] ^ codeword[863] ^ codeword[879] ^ codeword[880] ^ codeword[881] ^ codeword[882] ^ codeword[883] ^ codeword[884] ^ codeword[891] ^ codeword[912] ^ codeword[913] ^ codeword[914] ^ codeword[915] ^ codeword[916] ^ codeword[917] ^ codeword[918] ^ codeword[919] ^ codeword[920] ^ codeword[921] ^ codeword[922] ^ codeword[923] ^ codeword[924] ^ codeword[925] ^ codeword[926] ^ codeword[942] ^ codeword[943] ^ codeword[944] ^ codeword[945] ^ codeword[946] ^ codeword[947] ^ codeword[963] ^ codeword[964] ^ codeword[965] ^ codeword[966] ^ codeword[967] ^ codeword[968] ^ codeword[975] ^ codeword[991] ^ codeword[992] ^ codeword[993] ^ codeword[994] ^ codeword[995] ^ codeword[996] ^ codeword[1003] ^ codeword[1010] ^ codeword[1012] ^ codeword[1014] ^ codeword[1015] ^ codeword[1016] ^ codeword[1017] ^ codeword[1018] ^ codeword[1019] ^ codeword[1021] ^ codeword[1022] ^ codeword[1023] ^ codeword[1029];
    assign syndrome[6] = codeword[10] ^ codeword[11] ^ codeword[12] ^ codeword[13] ^ codeword[14] ^ codeword[15] ^ codeword[16] ^ codeword[17] ^ codeword[18] ^ codeword[19] ^ codeword[30] ^ codeword[31] ^ codeword[32] ^ codeword[33] ^ codeword[34] ^ codeword[45] ^ codeword[46] ^ codeword[47] ^ codeword[48] ^ codeword[49] ^ codeword[55] ^ codeword[66] ^ codeword[67] ^ codeword[68] ^ codeword[69] ^ codeword[70] ^ codeword[76] ^ codeword[82] ^ codeword[94] ^ codeword[95] ^ codeword[96] ^ codeword[97] ^ codeword[98] ^ codeword[104] ^ codeword[110] ^ codeword[117] ^ codeword[130] ^ codeword[131] ^ codeword[132] ^ codeword[133] ^ codeword[134] ^ codeword[140] ^ codeword[146] ^ codeword[153] ^ codeword[161] ^ codeword[175] ^ codeword[176] ^ codeword[177] ^ codeword[178] ^ codeword[179] ^ codeword[185] ^ codeword[191] ^ codeword[198] ^ codeword[206] ^ codeword[215] ^ codeword[221] ^ codeword[222] ^ codeword[223] ^ codeword[224] ^ codeword[225] ^ codeword[231] ^ codeword[232] ^ codeword[233] ^ codeword[234] ^ codeword[235] ^ codeword[236] ^ codeword[237] ^ codeword[238] ^ codeword[239] ^ codeword[240] ^ codeword[246] ^ codeword[247] ^ codeword[248] ^ codeword[249] ^ codeword[250] ^ codeword[251] ^ codeword[252] ^ codeword[253] ^ codeword[254] ^ codeword[255] ^ codeword[266] ^ codeword[267] ^ codeword[268] ^ codeword[269] ^ codeword[270] ^ codeword[271] ^ codeword[272] ^ codeword[273] ^ codeword[274] ^ codeword[275] ^ codeword[281] ^ codeword[282] ^ codeword[283] ^ codeword[284] ^ codeword[285] ^ codeword[286] ^ codeword[287] ^ codeword[288] ^ codeword[289] ^ codeword[290] ^ codeword[301] ^ codeword[302] ^ codeword[303] ^ codeword[304] ^ codeword[305] ^ codeword[306] ^ codeword[307] ^ codeword[308] ^ codeword[309] ^ codeword[310] ^ codeword[321] ^ codeword[322] ^ codeword[323] ^ codeword[324] ^ codeword[325] ^ codeword[326] ^ codeword[327] ^ codeword[328] ^ codeword[329] ^ codeword[330] ^ codeword[341] ^ codeword[342] ^ codeword[343] ^ codeword[344] ^ codeword[345] ^ codeword[351] ^ codeword[352] ^ codeword[353] ^ codeword[354] ^ codeword[355] ^ codeword[356] ^ codeword[357] ^ codeword[358] ^ codeword[359] ^ codeword[360] ^ codeword[371] ^ codeword[372] ^ codeword[373] ^ codeword[374] ^ codeword[375] ^ codeword[376] ^ codeword[377] ^ codeword[378] ^ codeword[379] ^ codeword[380] ^ codeword[391] ^ codeword[392] ^ codeword[393] ^ codeword[394] ^ codeword[395] ^ codeword[396] ^ codeword[397] ^ codeword[398] ^ codeword[399] ^ codeword[400] ^ codeword[411] ^ codeword[412] ^ codeword[413] ^ codeword[414] ^ codeword[415] ^ codeword[426] ^ codeword[427] ^ codeword[428] ^ codeword[429] ^ codeword[430] ^ codeword[431] ^ codeword[432] ^ codeword[433] ^ codeword[434] ^ codeword[435] ^ codeword[446] ^ codeword[447] ^ codeword[448] ^ codeword[449] ^ codeword[450] ^ codeword[461] ^ codeword[462] ^ codeword[463] ^ codeword[464] ^ codeword[465] ^ codeword[471] ^ codeword[477] ^ codeword[478] ^ codeword[479] ^ codeword[480] ^ codeword[481] ^ codeword[482] ^ codeword[483] ^ codeword[484] ^ codeword[485] ^ codeword[486] ^ codeword[497] ^ codeword[498] ^ codeword[499] ^ codeword[500] ^ codeword[501] ^ codeword[502] ^ codeword[503] ^ codeword[504] ^ codeword[505] ^ codeword[506] ^ codeword[517] ^ codeword[518] ^ codeword[519] ^ codeword[520] ^ codeword[521] ^ codeword[522] ^ codeword[523] ^ codeword[524] ^ codeword[525] ^ codeword[526] ^ codeword[537] ^ codeword[538] ^ codeword[539] ^ codeword[540] ^ codeword[541] ^ codeword[552] ^ codeword[553] ^ codeword[554] ^ codeword[555] ^ codeword[556] ^ codeword[557] ^ codeword[558] ^ codeword[559] ^ codeword[560] ^ codeword[561] ^ codeword[572] ^ codeword[573] ^ codeword[574] ^ codeword[575] ^ codeword[576] ^ codeword[587] ^ codeword[588] ^ codeword[589] ^ codeword[590] ^ codeword[591] ^ codeword[597] ^ codeword[608] ^ codeword[609] ^ codeword[610] ^ codeword[611] ^ codeword[612] ^ codeword[613] ^ codeword[614] ^ codeword[615] ^ codeword[616] ^ codeword[617] ^ codeword[628] ^ codeword[629] ^ codeword[630] ^ codeword[631] ^ codeword[632] ^ codeword[643] ^ codeword[644] ^ codeword[645] ^ codeword[646] ^ codeword[647] ^ codeword[653] ^ codeword[664] ^ codeword[665] ^ codeword[666] ^ codeword[667] ^ codeword[668] ^ codeword[674] ^ codeword[680] ^ codeword[687] ^ codeword[688] ^ codeword[689] ^ codeword[690] ^ codeword[691] ^ codeword[692] ^ codeword[693] ^ codeword[694] ^ codeword[695] ^ codeword[696] ^ codeword[707] ^ codeword[708] ^ codeword[709] ^ codeword[710] ^ codeword[711] ^ codeword[712] ^ codeword[713] ^ codeword[714] ^ codeword[715] ^ codeword[716] ^ codeword[727] ^ codeword[728] ^ codeword[729] ^ codeword[730] ^ codeword[731] ^ codeword[732] ^ codeword[733] ^ codeword[734] ^ codeword[735] ^ codeword[736] ^ codeword[747] ^ codeword[748] ^ codeword[749] ^ codeword[750] ^ codeword[751] ^ codeword[762] ^ codeword[763] ^ codeword[764] ^ codeword[765] ^ codeword[766] ^ codeword[767] ^ codeword[768] ^ codeword[769] ^ codeword[770] ^ codeword[771] ^ codeword[782] ^ codeword[783] ^ codeword[784] ^ codeword[785] ^ codeword[786] ^ codeword[797] ^ codeword[798] ^ codeword[799] ^ codeword[800] ^ codeword[801] ^ codeword[807] ^ codeword[818] ^ codeword[819] ^ codeword[820] ^ codeword[821] ^ codeword[822] ^ codeword[823] ^ codeword[824] ^ codeword[825] ^ codeword[826] ^ codeword[827] ^ codeword[838] ^ codeword[839] ^ codeword[840] ^ codeword[841] ^ codeword[842] ^ codeword[853] ^ codeword[854] ^ codeword[855] ^ codeword[856] ^ codeword[857] ^ codeword[863] ^ codeword[874] ^ codeword[875] ^ codeword[876] ^ codeword[877] ^ codeword[878] ^ codeword[884] ^ codeword[890] ^ codeword[902] ^ codeword[903] ^ codeword[904] ^ codeword[905] ^ codeword[906] ^ codeword[907] ^ codeword[908] ^ codeword[909] ^ codeword[910] ^ codeword[911] ^ codeword[922] ^ codeword[923] ^ codeword[924] ^ codeword[925] ^ codeword[926] ^ codeword[937] ^ codeword[938] ^ codeword[939] ^ codeword[940] ^ codeword[941] ^ codeword[947] ^ codeword[958] ^ codeword[959] ^ codeword[960] ^ codeword[961] ^ codeword[962] ^ codeword[968] ^ codeword[974] ^ codeword[986] ^ codeword[987] ^ codeword[988] ^ codeword[989] ^ codeword[990] ^ codeword[996] ^ codeword[1002] ^ codeword[1009] ^ codeword[1012] ^ codeword[1013] ^ codeword[1015] ^ codeword[1016] ^ codeword[1017] ^ codeword[1018] ^ codeword[1019] ^ codeword[1020] ^ codeword[1022] ^ codeword[1023] ^ codeword[1030];
    assign syndrome[7] = codeword[4] ^ codeword[5] ^ codeword[6] ^ codeword[7] ^ codeword[8] ^ codeword[9] ^ codeword[16] ^ codeword[17] ^ codeword[18] ^ codeword[19] ^ codeword[26] ^ codeword[27] ^ codeword[28] ^ codeword[29] ^ codeword[34] ^ codeword[41] ^ codeword[42] ^ codeword[43] ^ codeword[44] ^ codeword[49] ^ codeword[54] ^ codeword[62] ^ codeword[63] ^ codeword[64] ^ codeword[65] ^ codeword[70] ^ codeword[75] ^ codeword[81] ^ codeword[90] ^ codeword[91] ^ codeword[92] ^ codeword[93] ^ codeword[98] ^ codeword[103] ^ codeword[109] ^ codeword[116] ^ codeword[126] ^ codeword[127] ^ codeword[128] ^ codeword[129] ^ codeword[134] ^ codeword[139] ^ codeword[145] ^ codeword[152] ^ codeword[160] ^ codeword[171] ^ codeword[172] ^ codeword[173] ^ codeword[174] ^ codeword[179] ^ codeword[184] ^ codeword[190] ^ codeword[197] ^ codeword[205] ^ codeword[214] ^ codeword[220] ^ codeword[222] ^ codeword[223] ^ codeword[224] ^ codeword[225] ^ codeword[227] ^ codeword[228] ^ codeword[229] ^ codeword[230] ^ codeword[235] ^ codeword[236] ^ codeword[237] ^ codeword[238] ^ codeword[239] ^ codeword[240] ^ codeword[242] ^ codeword[243] ^ codeword[244] ^ codeword[245] ^ codeword[250] ^ codeword[251] ^ codeword[252] ^ codeword[253] ^ codeword[254] ^ codeword[255] ^ codeword[260] ^ codeword[261] ^ codeword[262] ^ codeword[263] ^ codeword[264] ^ codeword[265] ^ codeword[272] ^ codeword[273] ^ codeword[274] ^ codeword[275] ^ codeword[277] ^ codeword[278] ^ codeword[279] ^ codeword[280] ^ codeword[285] ^ codeword[286] ^ codeword[287] ^ codeword[288] ^ codeword[289] ^ codeword[290] ^ codeword[295] ^ codeword[296] ^ codeword[297] ^ codeword[298] ^ codeword[299] ^ codeword[300] ^ codeword[307] ^ codeword[308] ^ codeword[309] ^ codeword[310] ^ codeword[315] ^ codeword[316] ^ codeword[317] ^ codeword[318] ^ codeword[319] ^ codeword[320] ^ codeword[327] ^ codeword[328] ^ codeword[329] ^ codeword[330] ^ codeword[337] ^ codeword[338] ^ codeword[339] ^ codeword[340] ^ codeword[345] ^ codeword[347] ^ codeword[348] ^ codeword[349] ^ codeword[350] ^ codeword[355] ^ codeword[356] ^ codeword[357] ^ codeword[358] ^ codeword[359] ^ codeword[360] ^ codeword[365] ^ codeword[366] ^ codeword[367] ^ codeword[368] ^ codeword[369] ^ codeword[370] ^ codeword[377] ^ codeword[378] ^ codeword[379] ^ codeword[380] ^ codeword[385] ^ codeword[386] ^ codeword[387] ^ codeword[388] ^ codeword[389] ^ codeword[390] ^ codeword[397] ^ codeword[398] ^ codeword[399] ^ codeword[400] ^ codeword[407] ^ codeword[408] ^ codeword[409] ^ codeword[410] ^ codeword[415] ^ codeword[420] ^ codeword[421] ^ codeword[422] ^ codeword[423] ^ codeword[424] ^ codeword[425] ^ codeword[432] ^ codeword[433] ^ codeword[434] ^ codeword[435] ^ codeword[442] ^ codeword[443] ^ codeword[444] ^ codeword[445] ^ codeword[450] ^ codeword[457] ^ codeword[458] ^ codeword[459] ^ codeword[460] ^ codeword[465] ^ codeword[470] ^ codeword[473] ^ codeword[474] ^ codeword[475] ^ codeword[476] ^ codeword[481] ^ codeword[482] ^ codeword[483] ^ codeword[484] ^ codeword[485] ^ codeword[486] ^ codeword[491] ^ codeword[492] ^ codeword[493] ^ codeword[494] ^ codeword[495] ^ codeword[496] ^ codeword[503] ^ codeword[504] ^ codeword[505] ^ codeword[506] ^ codeword[511] ^ codeword[512] ^ codeword[513] ^ codeword[514] ^ codeword[515] ^ codeword[516] ^ codeword[523] ^ codeword[524] ^ codeword[525] ^ codeword[526] ^ codeword[533] ^ codeword[534] ^ codeword[535] ^ codeword[536] ^ codeword[541] ^ codeword[546] ^ codeword[547] ^ codeword[548] ^ codeword[549] ^ codeword[550] ^ codeword[551] ^ codeword[558] ^ codeword[559] ^ codeword[560] ^ codeword[561] ^ codeword[568] ^ codeword[569] ^ codeword[570] ^ codeword[571] ^ codeword[576] ^ codeword[583] ^ codeword[584] ^ codeword[585] ^ codeword[586] ^ codeword[591] ^ codeword[596] ^ codeword[602] ^ codeword[603] ^ codeword[604] ^ codeword[605] ^ codeword[606] ^ codeword[607] ^ codeword[614] ^ codeword[615] ^ codeword[616] ^ codeword[617] ^ codeword[624] ^ codeword[625] ^ codeword[626] ^ codeword[627] ^ codeword[632] ^ codeword[639] ^ codeword[640] ^ codeword[641] ^ codeword[642] ^ codeword[647] ^ codeword[652] ^ codeword[660] ^ codeword[661] ^ codeword[662] ^ codeword[663] ^ codeword[668] ^ codeword[673] ^ codeword[679] ^ codeword[683] ^ codeword[684] ^ codeword[685] ^ codeword[686] ^ codeword[691] ^ codeword[692] ^ codeword[693] ^ codeword[694] ^ codeword[695] ^ codeword[696] ^ codeword[701] ^ codeword[702] ^ codeword[703] ^ codeword[704] ^ codeword[705] ^ codeword[706] ^ codeword[713] ^ codeword[714] ^ codeword[715] ^ codeword[716] ^ codeword[721] ^ codeword[722] ^ codeword[723] ^ codeword[724] ^ codeword[725] ^ codeword[726] ^ codeword[733] ^ codeword[734] ^ codeword[735] ^ codeword[736] ^ codeword[743] ^ codeword[744] ^ codeword[745] ^ codeword[746] ^ codeword[751] ^ codeword[756] ^ codeword[757] ^ codeword[758] ^ codeword[759] ^ codeword[760] ^ codeword[761] ^ codeword[768] ^ codeword[769] ^ codeword[770] ^ codeword[771] ^ codeword[778] ^ codeword[779] ^ codeword[780] ^ codeword[781] ^ codeword[786] ^ codeword[793] ^ codeword[794] ^ codeword[795] ^ codeword[796] ^ codeword[801] ^ codeword[806] ^ codeword[812] ^ codeword[813] ^ codeword[814] ^ codeword[815] ^ codeword[816] ^ codeword[817] ^ codeword[824] ^ codeword[825] ^ codeword[826] ^ codeword[827] ^ codeword[834] ^ codeword[835] ^ codeword[836] ^ codeword[837] ^ codeword[842] ^ codeword[849] ^ codeword[850] ^ codeword[851] ^ codeword[852] ^ codeword[857] ^ codeword[862] ^ codeword[870] ^ codeword[871] ^ codeword[872] ^ codeword[873] ^ codeword[878] ^ codeword[883] ^ codeword[889] ^ codeword[896] ^ codeword[897] ^ codeword[898] ^ codeword[899] ^ codeword[900] ^ codeword[901] ^ codeword[908] ^ codeword[909] ^ codeword[910] ^ codeword[911] ^ codeword[918] ^ codeword[919] ^ codeword[920] ^ codeword[921] ^ codeword[926] ^ codeword[933] ^ codeword[934] ^ codeword[935] ^ codeword[936] ^ codeword[941] ^ codeword[946] ^ codeword[954] ^ codeword[955] ^ codeword[956] ^ codeword[957] ^ codeword[962] ^ codeword[967] ^ codeword[973] ^ codeword[982] ^ codeword[983] ^ codeword[984] ^ codeword[985] ^ codeword[990] ^ codeword[995] ^ codeword[1001] ^ codeword[1008] ^ codeword[1012] ^ codeword[1013] ^ codeword[1014] ^ codeword[1016] ^ codeword[1017] ^ codeword[1018] ^ codeword[1019] ^ codeword[1020] ^ codeword[1021] ^ codeword[1023] ^ codeword[1031];
    assign syndrome[8] = codeword[1] ^ codeword[2] ^ codeword[3] ^ codeword[7] ^ codeword[8] ^ codeword[9] ^ codeword[13] ^ codeword[14] ^ codeword[15] ^ codeword[19] ^ codeword[23] ^ codeword[24] ^ codeword[25] ^ codeword[29] ^ codeword[33] ^ codeword[38] ^ codeword[39] ^ codeword[40] ^ codeword[44] ^ codeword[48] ^ codeword[53] ^ codeword[59] ^ codeword[60] ^ codeword[61] ^ codeword[65] ^ codeword[69] ^ codeword[74] ^ codeword[80] ^ codeword[87] ^ codeword[88] ^ codeword[89] ^ codeword[93] ^ codeword[97] ^ codeword[102] ^ codeword[108] ^ codeword[115] ^ codeword[123] ^ codeword[124] ^ codeword[125] ^ codeword[129] ^ codeword[133] ^ codeword[138] ^ codeword[144] ^ codeword[151] ^ codeword[159] ^ codeword[168] ^ codeword[169] ^ codeword[170] ^ codeword[174] ^ codeword[178] ^ codeword[183] ^ codeword[189] ^ codeword[196] ^ codeword[204] ^ codeword[213] ^ codeword[220] ^ codeword[221] ^ codeword[223] ^ codeword[224] ^ codeword[225] ^ codeword[226] ^ codeword[228] ^ codeword[229] ^ codeword[230] ^ codeword[232] ^ codeword[233] ^ codeword[234] ^ codeword[238] ^ codeword[239] ^ codeword[240] ^ codeword[241] ^ codeword[243] ^ codeword[244] ^ codeword[245] ^ codeword[247] ^ codeword[248] ^ codeword[249] ^ codeword[253] ^ codeword[254] ^ codeword[255] ^ codeword[257] ^ codeword[258] ^ codeword[259] ^ codeword[263] ^ codeword[264] ^ codeword[265] ^ codeword[269] ^ codeword[270] ^ codeword[271] ^ codeword[275] ^ codeword[276] ^ codeword[278] ^ codeword[279] ^ codeword[280] ^ codeword[282] ^ codeword[283] ^ codeword[284] ^ codeword[288] ^ codeword[289] ^ codeword[290] ^ codeword[292] ^ codeword[293] ^ codeword[294] ^ codeword[298] ^ codeword[299] ^ codeword[300] ^ codeword[304] ^ codeword[305] ^ codeword[306] ^ codeword[310] ^ codeword[312] ^ codeword[313] ^ codeword[314] ^ codeword[318] ^ codeword[319] ^ codeword[320] ^ codeword[324] ^ codeword[325] ^ codeword[326] ^ codeword[330] ^ codeword[334] ^ codeword[335] ^ codeword[336] ^ codeword[340] ^ codeword[344] ^ codeword[346] ^ codeword[348] ^ codeword[349] ^ codeword[350] ^ codeword[352] ^ codeword[353] ^ codeword[354] ^ codeword[358] ^ codeword[359] ^ codeword[360] ^ codeword[362] ^ codeword[363] ^ codeword[364] ^ codeword[368] ^ codeword[369] ^ codeword[370] ^ codeword[374] ^ codeword[375] ^ codeword[376] ^ codeword[380] ^ codeword[382] ^ codeword[383] ^ codeword[384] ^ codeword[388] ^ codeword[389] ^ codeword[390] ^ codeword[394] ^ codeword[395] ^ codeword[396] ^ codeword[400] ^ codeword[404] ^ codeword[405] ^ codeword[406] ^ codeword[410] ^ codeword[414] ^ codeword[417] ^ codeword[418] ^ codeword[419] ^ codeword[423] ^ codeword[424] ^ codeword[425] ^ codeword[429] ^ codeword[430] ^ codeword[431] ^ codeword[435] ^ codeword[439] ^ codeword[440] ^ codeword[441] ^ codeword[445] ^ codeword[449] ^ codeword[454] ^ codeword[455] ^ codeword[456] ^ codeword[460] ^ codeword[464] ^ codeword[469] ^ codeword[472] ^ codeword[474] ^ codeword[475] ^ codeword[476] ^ codeword[478] ^ codeword[479] ^ codeword[480] ^ codeword[484] ^ codeword[485] ^ codeword[486] ^ codeword[488] ^ codeword[489] ^ codeword[490] ^ codeword[494] ^ codeword[495] ^ codeword[496] ^ codeword[500] ^ codeword[501] ^ codeword[502] ^ codeword[506] ^ codeword[508] ^ codeword[509] ^ codeword[510] ^ codeword[514] ^ codeword[515] ^ codeword[516] ^ codeword[520] ^ codeword[521] ^ codeword[522] ^ codeword[526] ^ codeword[530] ^ codeword[531] ^ codeword[532] ^ codeword[536] ^ codeword[540] ^ codeword[543] ^ codeword[544] ^ codeword[545] ^ codeword[549] ^ codeword[550] ^ codeword[551] ^ codeword[555] ^ codeword[556] ^ codeword[557] ^ codeword[561] ^ codeword[565] ^ codeword[566] ^ codeword[567] ^ codeword[571] ^ codeword[575] ^ codeword[580] ^ codeword[581] ^ codeword[582] ^ codeword[586] ^ codeword[590] ^ codeword[595] ^ codeword[599] ^ codeword[600] ^ codeword[601] ^ codeword[605] ^ codeword[606] ^ codeword[607] ^ codeword[611] ^ codeword[612] ^ codeword[613] ^ codeword[617] ^ codeword[621] ^ codeword[622] ^ codeword[623] ^ codeword[627] ^ codeword[631] ^ codeword[636] ^ codeword[637] ^ codeword[638] ^ codeword[642] ^ codeword[646] ^ codeword[651] ^ codeword[657] ^ codeword[658] ^ codeword[659] ^ codeword[663] ^ codeword[667] ^ codeword[672] ^ codeword[678] ^ codeword[682] ^ codeword[684] ^ codeword[685] ^ codeword[686] ^ codeword[688] ^ codeword[689] ^ codeword[690] ^ codeword[694] ^ codeword[695] ^ codeword[696] ^ codeword[698] ^ codeword[699] ^ codeword[700] ^ codeword[704] ^ codeword[705] ^ codeword[706] ^ codeword[710] ^ codeword[711] ^ codeword[712] ^ codeword[716] ^ codeword[718] ^ codeword[719] ^ codeword[720] ^ codeword[724] ^ codeword[725] ^ codeword[726] ^ codeword[730] ^ codeword[731] ^ codeword[732] ^ codeword[736] ^ codeword[740] ^ codeword[741] ^ codeword[742] ^ codeword[746] ^ codeword[750] ^ codeword[753] ^ codeword[754] ^ codeword[755] ^ codeword[759] ^ codeword[760] ^ codeword[761] ^ codeword[765] ^ codeword[766] ^ codeword[767] ^ codeword[771] ^ codeword[775] ^ codeword[776] ^ codeword[777] ^ codeword[781] ^ codeword[785] ^ codeword[790] ^ codeword[791] ^ codeword[792] ^ codeword[796] ^ codeword[800] ^ codeword[805] ^ codeword[809] ^ codeword[810] ^ codeword[811] ^ codeword[815] ^ codeword[816] ^ codeword[817] ^ codeword[821] ^ codeword[822] ^ codeword[823] ^ codeword[827] ^ codeword[831] ^ codeword[832] ^ codeword[833] ^ codeword[837] ^ codeword[841] ^ codeword[846] ^ codeword[847] ^ codeword[848] ^ codeword[852] ^ codeword[856] ^ codeword[861] ^ codeword[867] ^ codeword[868] ^ codeword[869] ^ codeword[873] ^ codeword[877] ^ codeword[882] ^ codeword[888] ^ codeword[893] ^ codeword[894] ^ codeword[895] ^ codeword[899] ^ codeword[900] ^ codeword[901] ^ codeword[905] ^ codeword[906] ^ codeword[907] ^ codeword[911] ^ codeword[915] ^ codeword[916] ^ codeword[917] ^ codeword[921] ^ codeword[925] ^ codeword[930] ^ codeword[931] ^ codeword[932] ^ codeword[936] ^ codeword[940] ^ codeword[945] ^ codeword[951] ^ codeword[952] ^ codeword[953] ^ codeword[957] ^ codeword[961] ^ codeword[966] ^ codeword[972] ^ codeword[979] ^ codeword[980] ^ codeword[981] ^ codeword[985] ^ codeword[989] ^ codeword[994] ^ codeword[1000] ^ codeword[1007] ^ codeword[1012] ^ codeword[1013] ^ codeword[1014] ^ codeword[1015] ^ codeword[1017] ^ codeword[1018] ^ codeword[1019] ^ codeword[1020] ^ codeword[1021] ^ codeword[1022] ^ codeword[1032];
    assign syndrome[9] = codeword[0] ^ codeword[2] ^ codeword[3] ^ codeword[5] ^ codeword[6] ^ codeword[9] ^ codeword[11] ^ codeword[12] ^ codeword[15] ^ codeword[18] ^ codeword[21] ^ codeword[22] ^ codeword[25] ^ codeword[28] ^ codeword[32] ^ codeword[36] ^ codeword[37] ^ codeword[40] ^ codeword[43] ^ codeword[47] ^ codeword[52] ^ codeword[57] ^ codeword[58] ^ codeword[61] ^ codeword[64] ^ codeword[68] ^ codeword[73] ^ codeword[79] ^ codeword[85] ^ codeword[86] ^ codeword[89] ^ codeword[92] ^ codeword[96] ^ codeword[101] ^ codeword[107] ^ codeword[114] ^ codeword[121] ^ codeword[122] ^ codeword[125] ^ codeword[128] ^ codeword[132] ^ codeword[137] ^ codeword[143] ^ codeword[150] ^ codeword[158] ^ codeword[166] ^ codeword[167] ^ codeword[170] ^ codeword[173] ^ codeword[177] ^ codeword[182] ^ codeword[188] ^ codeword[195] ^ codeword[203] ^ codeword[212] ^ codeword[220] ^ codeword[221] ^ codeword[222] ^ codeword[224] ^ codeword[225] ^ codeword[226] ^ codeword[227] ^ codeword[229] ^ codeword[230] ^ codeword[231] ^ codeword[233] ^ codeword[234] ^ codeword[236] ^ codeword[237] ^ codeword[240] ^ codeword[241] ^ codeword[242] ^ codeword[244] ^ codeword[245] ^ codeword[246] ^ codeword[248] ^ codeword[249] ^ codeword[251] ^ codeword[252] ^ codeword[255] ^ codeword[256] ^ codeword[258] ^ codeword[259] ^ codeword[261] ^ codeword[262] ^ codeword[265] ^ codeword[267] ^ codeword[268] ^ codeword[271] ^ codeword[274] ^ codeword[276] ^ codeword[277] ^ codeword[279] ^ codeword[280] ^ codeword[281] ^ codeword[283] ^ codeword[284] ^ codeword[286] ^ codeword[287] ^ codeword[290] ^ codeword[291] ^ codeword[293] ^ codeword[294] ^ codeword[296] ^ codeword[297] ^ codeword[300] ^ codeword[302] ^ codeword[303] ^ codeword[306] ^ codeword[309] ^ codeword[311] ^ codeword[313] ^ codeword[314] ^ codeword[316] ^ codeword[317] ^ codeword[320] ^ codeword[322] ^ codeword[323] ^ codeword[326] ^ codeword[329] ^ codeword[332] ^ codeword[333] ^ codeword[336] ^ codeword[339] ^ codeword[343] ^ codeword[346] ^ codeword[347] ^ codeword[349] ^ codeword[350] ^ codeword[351] ^ codeword[353] ^ codeword[354] ^ codeword[356] ^ codeword[357] ^ codeword[360] ^ codeword[361] ^ codeword[363] ^ codeword[364] ^ codeword[366] ^ codeword[367] ^ codeword[370] ^ codeword[372] ^ codeword[373] ^ codeword[376] ^ codeword[379] ^ codeword[381] ^ codeword[383] ^ codeword[384] ^ codeword[386] ^ codeword[387] ^ codeword[390] ^ codeword[392] ^ codeword[393] ^ codeword[396] ^ codeword[399] ^ codeword[402] ^ codeword[403] ^ codeword[406] ^ codeword[409] ^ codeword[413] ^ codeword[416] ^ codeword[418] ^ codeword[419] ^ codeword[421] ^ codeword[422] ^ codeword[425] ^ codeword[427] ^ codeword[428] ^ codeword[431] ^ codeword[434] ^ codeword[437] ^ codeword[438] ^ codeword[441] ^ codeword[444] ^ codeword[448] ^ codeword[452] ^ codeword[453] ^ codeword[456] ^ codeword[459] ^ codeword[463] ^ codeword[468] ^ codeword[472] ^ codeword[473] ^ codeword[475] ^ codeword[476] ^ codeword[477] ^ codeword[479] ^ codeword[480] ^ codeword[482] ^ codeword[483] ^ codeword[486] ^ codeword[487] ^ codeword[489] ^ codeword[490] ^ codeword[492] ^ codeword[493] ^ codeword[496] ^ codeword[498] ^ codeword[499] ^ codeword[502] ^ codeword[505] ^ codeword[507] ^ codeword[509] ^ codeword[510] ^ codeword[512] ^ codeword[513] ^ codeword[516] ^ codeword[518] ^ codeword[519] ^ codeword[522] ^ codeword[525] ^ codeword[528] ^ codeword[529] ^ codeword[532] ^ codeword[535] ^ codeword[539] ^ codeword[542] ^ codeword[544] ^ codeword[545] ^ codeword[547] ^ codeword[548] ^ codeword[551] ^ codeword[553] ^ codeword[554] ^ codeword[557] ^ codeword[560] ^ codeword[563] ^ codeword[564] ^ codeword[567] ^ codeword[570] ^ codeword[574] ^ codeword[578] ^ codeword[579] ^ codeword[582] ^ codeword[585] ^ codeword[589] ^ codeword[594] ^ codeword[598] ^ codeword[600] ^ codeword[601] ^ codeword[603] ^ codeword[604] ^ codeword[607] ^ codeword[609] ^ codeword[610] ^ codeword[613] ^ codeword[616] ^ codeword[619] ^ codeword[620] ^ codeword[623] ^ codeword[626] ^ codeword[630] ^ codeword[634] ^ codeword[635] ^ codeword[638] ^ codeword[641] ^ codeword[645] ^ codeword[650] ^ codeword[655] ^ codeword[656] ^ codeword[659] ^ codeword[662] ^ codeword[666] ^ codeword[671] ^ codeword[677] ^ codeword[682] ^ codeword[683] ^ codeword[685] ^ codeword[686] ^ codeword[687] ^ codeword[689] ^ codeword[690] ^ codeword[692] ^ codeword[693] ^ codeword[696] ^ codeword[697] ^ codeword[699] ^ codeword[700] ^ codeword[702] ^ codeword[703] ^ codeword[706] ^ codeword[708] ^ codeword[709] ^ codeword[712] ^ codeword[715] ^ codeword[717] ^ codeword[719] ^ codeword[720] ^ codeword[722] ^ codeword[723] ^ codeword[726] ^ codeword[728] ^ codeword[729] ^ codeword[732] ^ codeword[735] ^ codeword[738] ^ codeword[739] ^ codeword[742] ^ codeword[745] ^ codeword[749] ^ codeword[752] ^ codeword[754] ^ codeword[755] ^ codeword[757] ^ codeword[758] ^ codeword[761] ^ codeword[763] ^ codeword[764] ^ codeword[767] ^ codeword[770] ^ codeword[773] ^ codeword[774] ^ codeword[777] ^ codeword[780] ^ codeword[784] ^ codeword[788] ^ codeword[789] ^ codeword[792] ^ codeword[795] ^ codeword[799] ^ codeword[804] ^ codeword[808] ^ codeword[810] ^ codeword[811] ^ codeword[813] ^ codeword[814] ^ codeword[817] ^ codeword[819] ^ codeword[820] ^ codeword[823] ^ codeword[826] ^ codeword[829] ^ codeword[830] ^ codeword[833] ^ codeword[836] ^ codeword[840] ^ codeword[844] ^ codeword[845] ^ codeword[848] ^ codeword[851] ^ codeword[855] ^ codeword[860] ^ codeword[865] ^ codeword[866] ^ codeword[869] ^ codeword[872] ^ codeword[876] ^ codeword[881] ^ codeword[887] ^ codeword[892] ^ codeword[894] ^ codeword[895] ^ codeword[897] ^ codeword[898] ^ codeword[901] ^ codeword[903] ^ codeword[904] ^ codeword[907] ^ codeword[910] ^ codeword[913] ^ codeword[914] ^ codeword[917] ^ codeword[920] ^ codeword[924] ^ codeword[928] ^ codeword[929] ^ codeword[932] ^ codeword[935] ^ codeword[939] ^ codeword[944] ^ codeword[949] ^ codeword[950] ^ codeword[953] ^ codeword[956] ^ codeword[960] ^ codeword[965] ^ codeword[971] ^ codeword[977] ^ codeword[978] ^ codeword[981] ^ codeword[984] ^ codeword[988] ^ codeword[993] ^ codeword[999] ^ codeword[1006] ^ codeword[1012] ^ codeword[1013] ^ codeword[1014] ^ codeword[1015] ^ codeword[1016] ^ codeword[1018] ^ codeword[1019] ^ codeword[1020] ^ codeword[1021] ^ codeword[1022] ^ codeword[1023] ^ codeword[1033];
    assign syndrome[10] = codeword[0] ^ codeword[1] ^ codeword[3] ^ codeword[4] ^ codeword[6] ^ codeword[8] ^ codeword[10] ^ codeword[12] ^ codeword[14] ^ codeword[17] ^ codeword[20] ^ codeword[22] ^ codeword[24] ^ codeword[27] ^ codeword[31] ^ codeword[35] ^ codeword[37] ^ codeword[39] ^ codeword[42] ^ codeword[46] ^ codeword[51] ^ codeword[56] ^ codeword[58] ^ codeword[60] ^ codeword[63] ^ codeword[67] ^ codeword[72] ^ codeword[78] ^ codeword[84] ^ codeword[86] ^ codeword[88] ^ codeword[91] ^ codeword[95] ^ codeword[100] ^ codeword[106] ^ codeword[113] ^ codeword[120] ^ codeword[122] ^ codeword[124] ^ codeword[127] ^ codeword[131] ^ codeword[136] ^ codeword[142] ^ codeword[149] ^ codeword[157] ^ codeword[165] ^ codeword[167] ^ codeword[169] ^ codeword[172] ^ codeword[176] ^ codeword[181] ^ codeword[187] ^ codeword[194] ^ codeword[202] ^ codeword[211] ^ codeword[220] ^ codeword[221] ^ codeword[222] ^ codeword[223] ^ codeword[225] ^ codeword[226] ^ codeword[227] ^ codeword[228] ^ codeword[230] ^ codeword[231] ^ codeword[232] ^ codeword[234] ^ codeword[235] ^ codeword[237] ^ codeword[239] ^ codeword[241] ^ codeword[242] ^ codeword[243] ^ codeword[245] ^ codeword[246] ^ codeword[247] ^ codeword[249] ^ codeword[250] ^ codeword[252] ^ codeword[254] ^ codeword[256] ^ codeword[257] ^ codeword[259] ^ codeword[260] ^ codeword[262] ^ codeword[264] ^ codeword[266] ^ codeword[268] ^ codeword[270] ^ codeword[273] ^ codeword[276] ^ codeword[277] ^ codeword[278] ^ codeword[280] ^ codeword[281] ^ codeword[282] ^ codeword[284] ^ codeword[285] ^ codeword[287] ^ codeword[289] ^ codeword[291] ^ codeword[292] ^ codeword[294] ^ codeword[295] ^ codeword[297] ^ codeword[299] ^ codeword[301] ^ codeword[303] ^ codeword[305] ^ codeword[308] ^ codeword[311] ^ codeword[312] ^ codeword[314] ^ codeword[315] ^ codeword[317] ^ codeword[319] ^ codeword[321] ^ codeword[323] ^ codeword[325] ^ codeword[328] ^ codeword[331] ^ codeword[333] ^ codeword[335] ^ codeword[338] ^ codeword[342] ^ codeword[346] ^ codeword[347] ^ codeword[348] ^ codeword[350] ^ codeword[351] ^ codeword[352] ^ codeword[354] ^ codeword[355] ^ codeword[357] ^ codeword[359] ^ codeword[361] ^ codeword[362] ^ codeword[364] ^ codeword[365] ^ codeword[367] ^ codeword[369] ^ codeword[371] ^ codeword[373] ^ codeword[375] ^ codeword[378] ^ codeword[381] ^ codeword[382] ^ codeword[384] ^ codeword[385] ^ codeword[387] ^ codeword[389] ^ codeword[391] ^ codeword[393] ^ codeword[395] ^ codeword[398] ^ codeword[401] ^ codeword[403] ^ codeword[405] ^ codeword[408] ^ codeword[412] ^ codeword[416] ^ codeword[417] ^ codeword[419] ^ codeword[420] ^ codeword[422] ^ codeword[424] ^ codeword[426] ^ codeword[428] ^ codeword[430] ^ codeword[433] ^ codeword[436] ^ codeword[438] ^ codeword[440] ^ codeword[443] ^ codeword[447] ^ codeword[451] ^ codeword[453] ^ codeword[455] ^ codeword[458] ^ codeword[462] ^ codeword[467] ^ codeword[472] ^ codeword[473] ^ codeword[474] ^ codeword[476] ^ codeword[477] ^ codeword[478] ^ codeword[480] ^ codeword[481] ^ codeword[483] ^ codeword[485] ^ codeword[487] ^ codeword[488] ^ codeword[490] ^ codeword[491] ^ codeword[493] ^ codeword[495] ^ codeword[497] ^ codeword[499] ^ codeword[501] ^ codeword[504] ^ codeword[507] ^ codeword[508] ^ codeword[510] ^ codeword[511] ^ codeword[513] ^ codeword[515] ^ codeword[517] ^ codeword[519] ^ codeword[521] ^ codeword[524] ^ codeword[527] ^ codeword[529] ^ codeword[531] ^ codeword[534] ^ codeword[538] ^ codeword[542] ^ codeword[543] ^ codeword[545] ^ codeword[546] ^ codeword[548] ^ codeword[550] ^ codeword[552] ^ codeword[554] ^ codeword[556] ^ codeword[559] ^ codeword[562] ^ codeword[564] ^ codeword[566] ^ codeword[569] ^ codeword[573] ^ codeword[577] ^ codeword[579] ^ codeword[581] ^ codeword[584] ^ codeword[588] ^ codeword[593] ^ codeword[598] ^ codeword[599] ^ codeword[601] ^ codeword[602] ^ codeword[604] ^ codeword[606] ^ codeword[608] ^ codeword[610] ^ codeword[612] ^ codeword[615] ^ codeword[618] ^ codeword[620] ^ codeword[622] ^ codeword[625] ^ codeword[629] ^ codeword[633] ^ codeword[635] ^ codeword[637] ^ codeword[640] ^ codeword[644] ^ codeword[649] ^ codeword[654] ^ codeword[656] ^ codeword[658] ^ codeword[661] ^ codeword[665] ^ codeword[670] ^ codeword[676] ^ codeword[682] ^ codeword[683] ^ codeword[684] ^ codeword[686] ^ codeword[687] ^ codeword[688] ^ codeword[690] ^ codeword[691] ^ codeword[693] ^ codeword[695] ^ codeword[697] ^ codeword[698] ^ codeword[700] ^ codeword[701] ^ codeword[703] ^ codeword[705] ^ codeword[707] ^ codeword[709] ^ codeword[711] ^ codeword[714] ^ codeword[717] ^ codeword[718] ^ codeword[720] ^ codeword[721] ^ codeword[723] ^ codeword[725] ^ codeword[727] ^ codeword[729] ^ codeword[731] ^ codeword[734] ^ codeword[737] ^ codeword[739] ^ codeword[741] ^ codeword[744] ^ codeword[748] ^ codeword[752] ^ codeword[753] ^ codeword[755] ^ codeword[756] ^ codeword[758] ^ codeword[760] ^ codeword[762] ^ codeword[764] ^ codeword[766] ^ codeword[769] ^ codeword[772] ^ codeword[774] ^ codeword[776] ^ codeword[779] ^ codeword[783] ^ codeword[787] ^ codeword[789] ^ codeword[791] ^ codeword[794] ^ codeword[798] ^ codeword[803] ^ codeword[808] ^ codeword[809] ^ codeword[811] ^ codeword[812] ^ codeword[814] ^ codeword[816] ^ codeword[818] ^ codeword[820] ^ codeword[822] ^ codeword[825] ^ codeword[828] ^ codeword[830] ^ codeword[832] ^ codeword[835] ^ codeword[839] ^ codeword[843] ^ codeword[845] ^ codeword[847] ^ codeword[850] ^ codeword[854] ^ codeword[859] ^ codeword[864] ^ codeword[866] ^ codeword[868] ^ codeword[871] ^ codeword[875] ^ codeword[880] ^ codeword[886] ^ codeword[892] ^ codeword[893] ^ codeword[895] ^ codeword[896] ^ codeword[898] ^ codeword[900] ^ codeword[902] ^ codeword[904] ^ codeword[906] ^ codeword[909] ^ codeword[912] ^ codeword[914] ^ codeword[916] ^ codeword[919] ^ codeword[923] ^ codeword[927] ^ codeword[929] ^ codeword[931] ^ codeword[934] ^ codeword[938] ^ codeword[943] ^ codeword[948] ^ codeword[950] ^ codeword[952] ^ codeword[955] ^ codeword[959] ^ codeword[964] ^ codeword[970] ^ codeword[976] ^ codeword[978] ^ codeword[980] ^ codeword[983] ^ codeword[987] ^ codeword[992] ^ codeword[998] ^ codeword[1005] ^ codeword[1012] ^ codeword[1013] ^ codeword[1014] ^ codeword[1015] ^ codeword[1016] ^ codeword[1017] ^ codeword[1019] ^ codeword[1020] ^ codeword[1021] ^ codeword[1022] ^ codeword[1023] ^ codeword[1034];
    assign syndrome[11] = codeword[0] ^ codeword[1] ^ codeword[2] ^ codeword[4] ^ codeword[5] ^ codeword[7] ^ codeword[10] ^ codeword[11] ^ codeword[13] ^ codeword[16] ^ codeword[20] ^ codeword[21] ^ codeword[23] ^ codeword[26] ^ codeword[30] ^ codeword[35] ^ codeword[36] ^ codeword[38] ^ codeword[41] ^ codeword[45] ^ codeword[50] ^ codeword[56] ^ codeword[57] ^ codeword[59] ^ codeword[62] ^ codeword[66] ^ codeword[71] ^ codeword[77] ^ codeword[84] ^ codeword[85] ^ codeword[87] ^ codeword[90] ^ codeword[94] ^ codeword[99] ^ codeword[105] ^ codeword[112] ^ codeword[120] ^ codeword[121] ^ codeword[123] ^ codeword[126] ^ codeword[130] ^ codeword[135] ^ codeword[141] ^ codeword[148] ^ codeword[156] ^ codeword[165] ^ codeword[166] ^ codeword[168] ^ codeword[171] ^ codeword[175] ^ codeword[180] ^ codeword[186] ^ codeword[193] ^ codeword[201] ^ codeword[210] ^ codeword[220] ^ codeword[221] ^ codeword[222] ^ codeword[223] ^ codeword[224] ^ codeword[226] ^ codeword[227] ^ codeword[228] ^ codeword[229] ^ codeword[231] ^ codeword[232] ^ codeword[233] ^ codeword[235] ^ codeword[236] ^ codeword[238] ^ codeword[241] ^ codeword[242] ^ codeword[243] ^ codeword[244] ^ codeword[246] ^ codeword[247] ^ codeword[248] ^ codeword[250] ^ codeword[251] ^ codeword[253] ^ codeword[256] ^ codeword[257] ^ codeword[258] ^ codeword[260] ^ codeword[261] ^ codeword[263] ^ codeword[266] ^ codeword[267] ^ codeword[269] ^ codeword[272] ^ codeword[276] ^ codeword[277] ^ codeword[278] ^ codeword[279] ^ codeword[281] ^ codeword[282] ^ codeword[283] ^ codeword[285] ^ codeword[286] ^ codeword[288] ^ codeword[291] ^ codeword[292] ^ codeword[293] ^ codeword[295] ^ codeword[296] ^ codeword[298] ^ codeword[301] ^ codeword[302] ^ codeword[304] ^ codeword[307] ^ codeword[311] ^ codeword[312] ^ codeword[313] ^ codeword[315] ^ codeword[316] ^ codeword[318] ^ codeword[321] ^ codeword[322] ^ codeword[324] ^ codeword[327] ^ codeword[331] ^ codeword[332] ^ codeword[334] ^ codeword[337] ^ codeword[341] ^ codeword[346] ^ codeword[347] ^ codeword[348] ^ codeword[349] ^ codeword[351] ^ codeword[352] ^ codeword[353] ^ codeword[355] ^ codeword[356] ^ codeword[358] ^ codeword[361] ^ codeword[362] ^ codeword[363] ^ codeword[365] ^ codeword[366] ^ codeword[368] ^ codeword[371] ^ codeword[372] ^ codeword[374] ^ codeword[377] ^ codeword[381] ^ codeword[382] ^ codeword[383] ^ codeword[385] ^ codeword[386] ^ codeword[388] ^ codeword[391] ^ codeword[392] ^ codeword[394] ^ codeword[397] ^ codeword[401] ^ codeword[402] ^ codeword[404] ^ codeword[407] ^ codeword[411] ^ codeword[416] ^ codeword[417] ^ codeword[418] ^ codeword[420] ^ codeword[421] ^ codeword[423] ^ codeword[426] ^ codeword[427] ^ codeword[429] ^ codeword[432] ^ codeword[436] ^ codeword[437] ^ codeword[439] ^ codeword[442] ^ codeword[446] ^ codeword[451] ^ codeword[452] ^ codeword[454] ^ codeword[457] ^ codeword[461] ^ codeword[466] ^ codeword[472] ^ codeword[473] ^ codeword[474] ^ codeword[475] ^ codeword[477] ^ codeword[478] ^ codeword[479] ^ codeword[481] ^ codeword[482] ^ codeword[484] ^ codeword[487] ^ codeword[488] ^ codeword[489] ^ codeword[491] ^ codeword[492] ^ codeword[494] ^ codeword[497] ^ codeword[498] ^ codeword[500] ^ codeword[503] ^ codeword[507] ^ codeword[508] ^ codeword[509] ^ codeword[511] ^ codeword[512] ^ codeword[514] ^ codeword[517] ^ codeword[518] ^ codeword[520] ^ codeword[523] ^ codeword[527] ^ codeword[528] ^ codeword[530] ^ codeword[533] ^ codeword[537] ^ codeword[542] ^ codeword[543] ^ codeword[544] ^ codeword[546] ^ codeword[547] ^ codeword[549] ^ codeword[552] ^ codeword[553] ^ codeword[555] ^ codeword[558] ^ codeword[562] ^ codeword[563] ^ codeword[565] ^ codeword[568] ^ codeword[572] ^ codeword[577] ^ codeword[578] ^ codeword[580] ^ codeword[583] ^ codeword[587] ^ codeword[592] ^ codeword[598] ^ codeword[599] ^ codeword[600] ^ codeword[602] ^ codeword[603] ^ codeword[605] ^ codeword[608] ^ codeword[609] ^ codeword[611] ^ codeword[614] ^ codeword[618] ^ codeword[619] ^ codeword[621] ^ codeword[624] ^ codeword[628] ^ codeword[633] ^ codeword[634] ^ codeword[636] ^ codeword[639] ^ codeword[643] ^ codeword[648] ^ codeword[654] ^ codeword[655] ^ codeword[657] ^ codeword[660] ^ codeword[664] ^ codeword[669] ^ codeword[675] ^ codeword[682] ^ codeword[683] ^ codeword[684] ^ codeword[685] ^ codeword[687] ^ codeword[688] ^ codeword[689] ^ codeword[691] ^ codeword[692] ^ codeword[694] ^ codeword[697] ^ codeword[698] ^ codeword[699] ^ codeword[701] ^ codeword[702] ^ codeword[704] ^ codeword[707] ^ codeword[708] ^ codeword[710] ^ codeword[713] ^ codeword[717] ^ codeword[718] ^ codeword[719] ^ codeword[721] ^ codeword[722] ^ codeword[724] ^ codeword[727] ^ codeword[728] ^ codeword[730] ^ codeword[733] ^ codeword[737] ^ codeword[738] ^ codeword[740] ^ codeword[743] ^ codeword[747] ^ codeword[752] ^ codeword[753] ^ codeword[754] ^ codeword[756] ^ codeword[757] ^ codeword[759] ^ codeword[762] ^ codeword[763] ^ codeword[765] ^ codeword[768] ^ codeword[772] ^ codeword[773] ^ codeword[775] ^ codeword[778] ^ codeword[782] ^ codeword[787] ^ codeword[788] ^ codeword[790] ^ codeword[793] ^ codeword[797] ^ codeword[802] ^ codeword[808] ^ codeword[809] ^ codeword[810] ^ codeword[812] ^ codeword[813] ^ codeword[815] ^ codeword[818] ^ codeword[819] ^ codeword[821] ^ codeword[824] ^ codeword[828] ^ codeword[829] ^ codeword[831] ^ codeword[834] ^ codeword[838] ^ codeword[843] ^ codeword[844] ^ codeword[846] ^ codeword[849] ^ codeword[853] ^ codeword[858] ^ codeword[864] ^ codeword[865] ^ codeword[867] ^ codeword[870] ^ codeword[874] ^ codeword[879] ^ codeword[885] ^ codeword[892] ^ codeword[893] ^ codeword[894] ^ codeword[896] ^ codeword[897] ^ codeword[899] ^ codeword[902] ^ codeword[903] ^ codeword[905] ^ codeword[908] ^ codeword[912] ^ codeword[913] ^ codeword[915] ^ codeword[918] ^ codeword[922] ^ codeword[927] ^ codeword[928] ^ codeword[930] ^ codeword[933] ^ codeword[937] ^ codeword[942] ^ codeword[948] ^ codeword[949] ^ codeword[951] ^ codeword[954] ^ codeword[958] ^ codeword[963] ^ codeword[969] ^ codeword[976] ^ codeword[977] ^ codeword[979] ^ codeword[982] ^ codeword[986] ^ codeword[991] ^ codeword[997] ^ codeword[1004] ^ codeword[1012] ^ codeword[1013] ^ codeword[1014] ^ codeword[1015] ^ codeword[1016] ^ codeword[1017] ^ codeword[1018] ^ codeword[1020] ^ codeword[1021] ^ codeword[1022] ^ codeword[1023] ^ codeword[1035];
  end else begin : gen_default_parity
    `BR_ASSERT_STATIC(invalid_parity_width_a, 1'b0)
  end
  // verilog_lint: waive-stop line-length
  // verilog_format: on


  // Decode syndrome.
  // * Case 0: Syndrome is zero, no errors detected.
  // * Case 1: Syndrome is for an even number of bits in error, which happens when the syndrome is even in a Hsiao SECDED code.
  //   Maximum likelihood decoding produces multiple equiprobable candidate codewords, so treat as detected-but-uncorrectable.
  //   NOTE: We are returning *some* message but it is likely to have been corrupted!
  // * Remaining case: Syndrome is for an odd number of bits in error, which happens when the syndrome is odd in a Hsiao SECDED code.
  //   *Usually* this is a single-bit error, which is always closest to exactly one codeword. So with maximum likelihood decoding
  //   we can correct it. However, sometimes it can be a three-bit error that is actually detected-but-uncorrectable.

  logic [ParityWidth-1:0] syndrome_ones_count;
  logic syndrome_is_zero;
  logic syndrome_is_even;
  logic syndrome_is_odd;
  logic [CodewordWidth-1:0] column_match_onehot;

  br_enc_countones #(
      .Width(ParityWidth)
  ) br_enc_countones_syndrome (
      .in(error_syndrome),
      .count(syndrome_ones_count)
  );

  assign syndrome_is_zero = error_syndrome == '0;
  assign syndrome_is_even = !syndrome_is_zero && !syndrome_ones_count[0];
  assign syndrome_is_odd = syndrome_ones_count[1];

  // TODO(mgottscho): Implement this. Need code generation. (WIP)
  assign column_match_onehot = '0;

  assign error_detected_but_uncorrectable = codeword_valid &&
    (syndrome_is_even || (syndrome_is_odd && column_match_onehot == 0));
  assign error_corrected = codeword_valid && syndrome_is_odd && (column_match_onehot != 0);

  // Actually correct the error.
  logic PadWidth = MessageWidth - DataWidth;
  logic [CodewordWidth-1:0] corrected_codeword;
  logic [MessageWidth-1:0] message;

  assign corrected_codeword = codeword ^ column_match_onehot;

  assign message = corrected_codeword[MessageWidth-1:0];
  assign data_valid = codeword_valid;
  assign data = message[DataWidth-1:0];

  //------------------------------------------
  // Implementation checks
  //------------------------------------------
  `BR_ASSERT_COMB_IMPL(data_valid_only_if_codeword_valid_a, !data_valid || codeword_valid)
  `BR_ASSERT_COMB_IMPL(error_valid_only_if_data_valid_a, !error_valid || data_valid)
  `BR_ASSERT_COMB_IMPL(ce_due_mutually_exclusive_a,
                       !error_valid || !(error_corrected && error_detected_but_uncorrectable))
  `BR_COVER_COMB_IMPL(error_valid_c, error_valid)
  `BR_COVER_COMB_IMPL(ce_c, error_valid && error_corrected)
  `BR_COVER_COMB_IMPL(due_c, error_valid && error_detected_but_uncorrectable)

endmodule : br_ecc_secded_decoder
