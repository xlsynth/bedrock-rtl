
// SPDX-License-Identifier: Apache-2.0
//
// Bedrock-RTL Shared Pseudo-Static Multi-FIFO w/ Flop-based Storage
// (Push Valid/Ready Interface, Pop Ready/Valid Interface)
//
// This module implements a shared storage multi-FIFO with flop-based storage.
// and pseudo-static allocation.
//
// The multi-FIFO contains multiple logical FIFOs. Space in the shared
// data RAM is allocated to the logical FIFOs statically at initialization,
// and a separate set of read/write pointers are kept per logical FIFO.
// For instance, for a 4-FIFO design with a depth of 16, the sizes of the
// logical FIFOs might be [6, 2, 3, 5]. In this case, you would configure
// the base and bound addresses as [(0, 5), (6, 7), (8, 10), (11, 15)] and the
// layout of the data RAM is as follows:
//
//  +----------------------------------------------------------------------------+
//  | Addr | 0 | 1 | 2 | 3 | 4 | 5 | 6 | 7 | 8 | 9 | 10 | 11 | 12 | 13 | 14 | 15 |
//  |------|---|---|---|---|---|---|---|---|---|---|----|----|----|----|----|----|
//  | FIFO | 0 | 0 | 0 | 0 | 0 | 0 | 1 | 1 | 2 | 2 | 2  | 3  | 3  | 3  | 3  | 3  |
//  +----------------------------------------------------------------------------+
//
// The push interface provides a valid/ready interface and a binary-encoded
// FIFO ID. The push data is appended to the logical FIFO with the specified ID.
//
//
// Every logical FIFO has its own ready/valid pop interface. If the data RAM
// read latency is non-zero or the RegisterPopOutputs parameter is set to 1, the
// pop_data will be provided from a staging buffer per logical FIFO. The staging
// buffers are refilled from the data RAM and arbitrate with each other for
// access. The depth of each staging buffer can be configured with the
// StagingBufferDepth parameter. The bandwidth of a single logical FIFO is
// determined by the staging buffer depth and is equivalent to
// `StagingBufferDepth / (RamReadLatency + 1)`.
//
// The design uses internal flop-based RAMs for the data storage.
// The latency of the internal RAM is determined from the retiming parameters as follows:
//
// `RamReadLatency = RamAddressDepthStages + RamReadDataDepthStages + RamReadDataWidthStages`
//
// The design uses internal arbiters to determine which logical FIFOs can use the RAM read ports
// on a given cycle. The arbitration policy is least-recently used (LRU).

`include "br_asserts_internal.svh"

// ri lint_check_waive MOD_NAME
module br_fifo_shared_pstatic_flops #(
    // Number of logical FIFOs. Must be >=2.
    parameter int NumFifos = 2,
    // Total depth of the FIFO.
    // Must be greater than two times the number of write ports.
    parameter int Depth = 2,
    // Width of the data. Must be >=1.
    parameter int Width = 1,
    // Number of write ports. Must be >=1.
    parameter int NumWritePorts = 1,
    // Number of read ports. Must be >=1 and a power of 2.
    parameter int NumReadPorts = 1,
    // The depth of the pop-side staging buffer.
    // This affects the pop bandwidth of each logical FIFO.
    // The max bandwidth will be `StagingBufferDepth / (DataRamReadLatency + 1)`.
    parameter int StagingBufferDepth = 1,
    // If 1, make sure pop_valid/pop_data are registered at the output
    // of the staging buffer. This adds a cycle of cut-through latency.
    parameter bit RegisterPopOutputs = 0,
    // If 1, place a register on the deallocation path from the pop-side
    // staging buffer to the freelist. This improves timing at the cost of
    // adding a cycle of backpressure latency.
    parameter bit RegisterDeallocation = 0,
    // Number of tiles in the depth dimension for the data flop RAM.
    parameter int RamDepthTiles = 1,
    // Number of tiles in the width dimension for the data flop RAM.
    parameter int RamWidthTiles = 1,
    // Number of stages on the address path for the data flop RAM.
    parameter int RamAddressDepthStages = 0,
    // Number of stages in the depth dimension on the data flop RAM.
    parameter int RamReadDataDepthStages = 0,
    // Number of stages in the width dimension on the data flop RAM.
    parameter int RamReadDataWidthStages = 0,
    // If 1, cover that the push side experiences backpressure.
    // If 0, assert that there is never backpressure.
    parameter bit EnableCoverPushBackpressure = 1,
    // If 1, assert that push_valid is stable when backpressured.
    parameter bit EnableAssertPushValidStability = EnableCoverPushBackpressure,
    // If 1, assert that push_data is stable when backpressured.
    // ri lint_check_waive PARAM_NOT_USED
    parameter bit EnableAssertPushDataStability = EnableAssertPushValidStability,
    // If 1, assert that push_data is always known (not X) when push_valid is asserted.
    parameter bit EnableAssertPushDataKnown = 1,
    // If 1, then assert there are no valid bits asserted and that the FIFO is
    // empty at the end of the test.
    // ri lint_check_waive PARAM_NOT_USED
    parameter bit EnableAssertFinalNotValid = 1,
    localparam int FifoIdWidth = br_math::clamped_clog2(NumFifos),
    localparam int AddrWidth = br_math::clamped_clog2(Depth)
) (
    input logic clk,
    input logic rst,
    // Fifo configuration
    // These can come from straps or CSRs, but they must be set before reset is
    // deasserted and then held stable until reset is asserted.
    // The base and bound addresses determine the range of RAM addresses given
    // to each logical FIFO. They are both inclusive, so logical FIFO i will
    // increment from config_base[i] up to config_bound[i] before wrapping back
    // around to config_base[i] again.
    // The minimum size for a given logical FIFO is 1, meaning that
    // config_bound[i] must be >= config_base[i] for all i.
    // The address ranges must be in ascending order.
    input logic [NumFifos-1:0][AddrWidth-1:0] config_base,
    input logic [NumFifos-1:0][AddrWidth-1:0] config_bound,
    // Error is asserted if the base and bound addresses are misconfigured.
    // For instance, if any address is >= Depth, config_base[i] > config_bound[i],
    // or config_base[i] <= config_bound[i-1] for i > 0.
    output logic config_error,

    // Push side
    output logic [NumWritePorts-1:0] push_ready,
    input logic [NumWritePorts-1:0] push_valid,
    input logic [NumWritePorts-1:0][Width-1:0] push_data,
    input logic [NumWritePorts-1:0][FifoIdWidth-1:0] push_fifo_id,
    output logic [NumFifos-1:0] push_full,

    // Pop side
    output logic [NumFifos-1:0] pop_valid,
    input logic [NumFifos-1:0] pop_ready,
    output logic [NumFifos-1:0][Width-1:0] pop_data,
    output logic [NumFifos-1:0] pop_empty
);

  // Integration Checks
  // Rely on checks in the submodules

  // Implementation
  // Data RAM
  logic ram_wr_valid;
  logic [AddrWidth-1:0] ram_wr_addr;
  logic [Width-1:0] ram_wr_data;

  logic ram_rd_addr_valid;
  logic [AddrWidth-1:0] ram_rd_addr;
  logic ram_rd_data_valid;
  logic [Width-1:0] ram_rd_data;

  br_ram_flops #(
      .Depth(Depth),
      .Width(Width),
      .NumWritePorts(1),
      .NumReadPorts(1),
      .DepthTiles(RamDepthTiles),
      .WidthTiles(RamWidthTiles),
      .AddressDepthStages(RamAddressDepthStages),
      .ReadDataDepthStages(RamReadDataDepthStages),
      .ReadDataWidthStages(RamReadDataWidthStages)
  ) br_ram_flops_data (
      .wr_clk(clk),  // ri lint_check_waive SAME_CLOCK_NAME
      .wr_rst(rst),
      .wr_valid(ram_wr_valid),
      .wr_addr(ram_wr_addr),
      .wr_data(ram_wr_data),
      .wr_word_en({RamWidthTiles{1'b1}}),
      .rd_clk(clk),  // ri lint_check_waive SAME_CLOCK_NAME
      .rd_rst(rst),
      .rd_addr_valid(ram_rd_addr_valid),
      .rd_addr(ram_rd_addr),
      .rd_data_valid(ram_rd_data_valid),
      .rd_data(ram_rd_data)
  );

  // Controller
  localparam int RamReadLatency =
      RamAddressDepthStages + RamReadDataDepthStages + RamReadDataWidthStages;

  br_fifo_shared_pstatic_ctrl #(
      .NumFifos(NumFifos),
      .Depth(Depth),
      .Width(Width),
      .NumWritePorts(NumWritePorts),
      .NumReadPorts(NumReadPorts),
      .StagingBufferDepth(StagingBufferDepth),
      .RegisterPopOutputs(RegisterPopOutputs),
      .RamReadLatency(RamReadLatency),
      .RegisterDeallocation(RegisterDeallocation),
      .EnableCoverPushBackpressure(EnableCoverPushBackpressure),
      .EnableAssertPushValidStability(EnableAssertPushValidStability),
      .EnableAssertPushDataStability(EnableAssertPushDataStability),
      .EnableAssertPushDataKnown(EnableAssertPushDataKnown),
      .EnableAssertFinalNotValid(EnableAssertFinalNotValid)
  ) br_fifo_shared_pstatic_ctrl_inst (
      .clk,
      .rst,
      .config_base,
      .config_bound,
      .config_error,
      .push_ready,
      .push_valid,
      .push_fifo_id,
      .push_data,
      .push_full,
      .pop_ready,
      .pop_valid,
      .pop_data,
      .pop_empty,
      .ram_wr_valid,
      .ram_wr_addr,
      .ram_wr_data,
      .ram_rd_addr_valid,
      .ram_rd_addr,
      .ram_rd_data_valid,
      .ram_rd_data
  );

  // Implementation Checks

  // Rely on implementation checks in the controller
endmodule : br_fifo_shared_pstatic_flops
